----------------------------------------------------------------------------------
-- Company: RIIC
-- Engineer: Gerhard Hohner Mat.nr.: 7555111
-- 
-- Create Date:    01/07/2004 
-- Design Name:    Diplomarbeit
-- Module Name:    ROMcode - Rtl 
-- Project Name:   32 bit FORTH processor
-- Target Devices: Spartan 3
-- Tool versions:  ISE 8.2
-- Description: implements a ROM containing the BIOS
-- Dependencies: global.vhd
-- 
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------


library IEEE, work;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.global.all;

entity ROMcode is
  port (Clock: in std_ulogic;									-- system clock
        Address: in std_ulogic_vector(ROMrange);		-- address bus
		  Data: out DataVec);									-- outgoing data
end ROMcode;

architecture RTL of ROMcode is
  type blocks is array (0 to 2048 / 4 - 1) of DataVec;
  type myarray is array (natural range <>) of blocks;
  constant ROM: myarray := (
(
"01000110010011100101011001010100",
"00001100001111100010010110000000",
"00000000000110110100011000100111",
"00000001111111111111000001000110",
"00111001000000000001011101000110",
"00000000000110000100011000000001",
"00001110010101100000000100110100",
"10010000000010100110010001000110",
"00011101100010000001000000000001",
"00000110001111100101001100000001",
"01000110000000100101101001000000",
"10000111001111100000001111101000",
"01000000010111010011111000010001",
"00000010111111111101010001000110",
"00000000000000000000110100001000",
"11011000000011010000011000000000",
"00000001000001011111111111111111",
"00001010010000000100011001010110",
"01000100010001100101011000000001",
"00001110010101100000000100001010",
"10010000000010100101100001000110",
"00011101100010000001000000000001",
"01111000010001100101011000000001",
"01000110010101100000000100001010",
"01010110000000010000101001111100",
"00000001010110101000100001000110",
"01011010100000000100011001001110",
"10000100010001100101011000000001",
"01000110010101100000000101011010",
"01000110000000010000101001100000",
"00001101010100100101101010010000",
"00000100000000000000110010001110",
"00000000000010111011100100111110",
"01010010010101100000000000000000",
"00000000000011001000100000001101",
"00001011101011000011111000000100",
"01001100000000000000000000000000",
"00001100100000100000110101010010",
"10011111001111100000010000000000",
"00000000000000000000000000001011",
"00000000000000000000000000001101",
"01111001000011010101001000000110",
"00111110000001000000000000001100",
"00000000000000000000101110001110",
"00000000000000000000110100000000",
"00001101010100100000011000000000",
"00000100000000000000110001101110",
"00000000000010110111110100111110",
"00010000010001100000000000000000",
"01100011000011010101001000000000",
"00111110000001000000000000001100",
"00000000000000000000101101101110",
"00001010011001000100011000000000",
"00001100010101010000110101010010",
"01011111001111100000010000000000",
"00000000000000000000000000001011",
"00000000000011000011110000001101",
"11000101000011010101001100000100",
"00111110000001000000000000001100",
"00010001000011010000101101001110",
"01010011000001000000000000001101",
"00000000000011010110001000001101",
"00001011010000000011111000000100",
"00000000000011010001110100001101",
"11000110000011010101001100000100",
"00111110000001000000000000001101",
"01101000000011010000101100110010",
"01010011000001000000000000001101",
"00000000000011100001011100001101",
"00001011001001000011111000000100",
"00000000000011100010000000001101",
"00101100000011010101001100000100",
"00111110000001000000000000001110",
"00100110000011010000101100010110",
"01010011000001000000000000001110",
"00000000000011100011101100001101",
"00001011000010000011111000000100",
"00000000000011100011011100001101",
"01101111000011010101001100000100",
"00111110000001000000000000001110",
"01000110000011010000101011111010",
"01010011000001000000000000001110",
"00000000000011100111100100001101",
"00001010111011000011111000000100",
"00000000000011100111010100001101",
"11110000000011010101001100000100",
"00111110000001000000000000001110",
"01001010000011010000101011011110",
"01010011000001000000000000001111",
"00000000000011111000100100001101",
"00001010110100000011111000000100",
"00000000000011111011111000001101",
"11011010000011010101001100000100",
"00111110000001000000000000001111",
"11001100000011010000101011000010",
"01010011000001000000000000001111",
"00000000000100000000000000001101",
"00001010101101000011111000000100",
"00000000000011111110000000001101",
"00001011000011010101001100000100",
"00111110000001000000000000010000",
"00000110000011010000101010100110",
"01010011000001000000000000010000",
"00000000000100000010011000001101",
"00001010100110000011111000000100",
"00000000000100000001001100001101",
"00111001000011010101001100000100",
"00111110000001000000000000010000",
"00101101000011010000101010001010",
"01010011000001000000000000010000",
"00000000000100001110001000001101",
"00001010011111000011111000000100",
"00000000000100000011110100001101",
"11111001000011010101001100000100",
"00111110000001000000000000010000",
"11101001000011010000101001101110",
"01010011000001000000000000010000",
"00000000000100010000011100001101",
"00001010011000000011111000000100",
"00000000000100010000001000001101",
"00110101000011010101001100000100",
"00111110000001000000000000010001",
"00001111000011010000101001010010",
"01010011000001000000000000010001",
"00000000000100010101001100001101",
"00001010010001000011111000000100",
"00000000000100010011110100001101",
"10011000000011010101001100000100",
"00111110000001000000000000010001",
"01011011000011010000101000110110",
"01010011000001000000000000010001",
"00000000000100011010010100001101",
"00001010001010000011111000000100",
"00000000000100011010000000001101",
"10110101000011010101001100000100",
"00111110000001000000000000010001",
"10101001000011010000101000011010",
"01010011000001000000000000010001",
"00000000000100011011110100001101",
"00001010000011000011111000000100",
"00000000000100011011100000001101",
"11001000000011010101001100000100",
"00111110000001000000000000010001",
"11000011000011010000100111111110",
"01010011000001000000000000010001",
"00000000000100011101011000001101",
"00001001111100000011111000000100",
"00000000000100011100101100001101",
"11100000000011010101001100000100",
"00111110000001000000000000010001",
"11011011000011010000100111100010",
"01010011000001000000000000010001",
"00000000000100101011010100001101",
"00001001110101000011111000000100",
"00000000000100011110011100001101",
"11001001000011010101001100000100",
"00111110000001000000000000010010",
"10111001000011010000100111000110",
"01010011000001000000000000010010",
"00000000000100110010010100001101",
"00001001101110000011111000000100",
"00000000000100101101001000001101",
"01110101000011010101001100000100",
"00111110000001000000000000010011",
"00101110000011010000100110101010",
"01010011000001000000000000010011",
"00000000000100111100001100001101",
"00001001100111000011111000000100",
"00000000000100110111110100001101",
"01000101000011010101001100000100",
"00111110000001000000000000010100",
"11001011000011010000100110001110",
"01010011000001000000000000010011",
"00000000000101001000101000001101",
"00001001100000000011111000000100",
"00000000000101000100110100001101",
"11000110000011010101001100000100",
"00111110000001000000000000010100",
"10001110000011010000100101110010",
"01010011000001000000000000010100",
"00000000000101001101010100001101",
"00001001011001000011111000000100",
"00000000000101001100101000001101",
"00011111000011010101001100000100",
"00111110000001000000000000010101",
"11011011000011010000100101010110",
"01010011000001000000000000010100",
"00000000000101010111100000001101",
"00001001010010000011111000000100",
"00000000000101010111110100001101",
"01001011000011010101001100000100",
"00111110000001000000000000010110",
"01010011000011010000100100111010",
"01010011000001000000000000010110",
"00000000000101110110000100001101",
"00001001001011000011111000000100",
"00000000000101111001011000001101",
"10001010000011010101001100000100",
"00111110000001000000000000011000",
"10000011000011010000100100011110",
"01010011000001000000000000011000",
"00000000000110100011001000001101",
"00001001000100000011111000000100",
"00000000000110001000111000001101",
"10011101000011010101001100000100",
"00111110000001000000000000011010",
"00110110000011010000100100000010",
"01010011000001000000000000011010",
"00000000000110110010011000001101",
"00001000111101000011111000000100",
"00000000000110101010000100001101",
"01110100000011010101001100000100",
"00111110000001000000000000011011",
"00110010000011010000100011100110",
"01010011000001000000000000011011",
"00000000000110111010000100001101",
"00001000110110000011111000000100",
"00000000000110110111100100001101",
"11001001000011010101001100000100",
"00111110000001000000000000011011",
"10101001000011010000100011001010",
"01010011000001000000000000011011",
"00000000000110111110111100001101",
"00001000101111000011111000000100",
"00000000000110111101000000001101",
"00011110000011010101001100000100",
"00111110000001000000000000011100",
"11110101000011010000100010101110",
"01010011000001000000000000011011",
"00000000000111000011010000001101",
"00001000101000000011111000000100",
"00000000000111000010010000001101",
"01010000000011010101001100000100",
"00111110000001000000000000011100",
"00111100000011010000100010010010",
"01010011000001000000000000011100",
"00000000000111000110111100001101",
"00001000100001000011111000000100",
"00000000000111000101010100001101",
"10000111000011010101001100000100",
"00111110000001000000000000011100",
"01110110000011010000100001110110",
"01010011000001000000000000011100",
"00000000000111001010110000001101",
"00001000011010000011111000000100",
"00000000000111001000111100001101",
"11001101000011010101001100000100",
"00111110000001000000000000011100",
"10110011000011010000100001011010",
"01010011000001000000000000011100",
"00000000000111010001111000001101",
"00001000010011000011111000000100",
"00000000000111001101010000001101",
"01001110000011010101001100000100",
"00111110000001000000000000011101",
"00100110000011010000100000111110",
"01010011000001000000000000011101",
"00000000000111010111110000001101",
"00001000001100000011111000000100",
"00000000000111010101010100001101",
"11001111000011010101001100000100",
"00111110000001000000000000011101",
"10000100000011010000100000100010",
"01010011000001000000000000011101",
"00000000000111011111010100001101",
"00001000000101000011111000000100",
"00000000000111011101011100001101",
"00111110000011010101001100000100",
"00111110000001000000000000011110",
"11111011000011010000100000000110",
"01010011000001000000000000011101",
"00000000000111100101001000001101",
"00000111111110000011111000000100",
"00000000000111100100010100001101",
"11110011000011010101001100000100",
"00111110000001000000000000011110",
"01011000000011010000011111101010",
"01010011000001000000000000011110",
"00000000000111110000100000001101",
"00000111110111000011111000000100",
"00000000000111101111101100001101",
"00011110000011010101001100000100",
"00111110000001000000000000011111",
"00001101000011010000011111001110",
"01010011000001000000000000011111",
"00000000000111110110111100001101",
"00000111110000000011111000000100",
"00000000000111110010010100001101",
"10010011000011010101001100000100",
"00111110000001000000000000011111",
"01110101000011010000011110110010",
"01010011000001000000000000011111",
"00000000000111111010010100001101",
"00000111101001000011111000000100",
"00000000000111111001100100001101",
"11111111000011010101001100000100",
"00111110000001000000000000011111",
"10101100000011010000011110010110",
"01010011000001000000000000011111",
"00000000001000000000111100001101",
"00000111100010000011111000000100",
"00000000001000000000100000001101",
"00111000000011010101001100000100",
"00111110000001000000000000100000",
"00010110000011010000011101111010",
"01010011000001000000000000100000",
"00000000001000000110011000001101",
"00000111011011000011111000000100",
"00000000001000000011111000001101",
"11001101000011010101001100000100",
"00111110000001000000000000100000",
"01101101000011010000011101011110",
"01010011000001000000000000100000",
"00000000001000001101100000001101",
"00000111010100000011111000000100",
"00000000001000001101000100001101",
"11111111000011010101001100000100",
"00111110000001000000000000100000",
"11011101000011010000011101000010",
"01010011000001000000000000100000",
"00000000001000010000101000001101",
"00000111001101000011111000000100",
"00000000001000010000001100001101",
"01000000000011010101001100000100",
"00111110000001000000000000100001",
"00010000000011010000011100100110",
"01010011000001000000000000100001",
"00000000001000010100110000001101",
"00000111000110000011111000000100",
"00000000001000010100010100001101",
"01110001000011010101001100000100",
"00111110000001000000000000100001",
"01010010000011010000011100001010",
"01010011000001000000000000100001",
"00000000001000011000100100001101",
"00000110111111000011111000000100",
"00000000001000111110110000001101",
"00000100000011010101001100000100",
"00111110000001000000000000100100",
"11111000000011010000011011101110",
"01010011000001000000000000100011",
"00000000001001000001001100001101",
"00000110111000000011111000000100",
"00000000001001000000100000001101",
"00111111000011010101001100000100",
"00111110000001000000000000100100",
"00011001000011010000011011010010",
"01010011000001000000000000100100",
"00000000001001000101000000001101",
"00000110110001000011111000000100",
"00000000001001000100010100001101",
"01100010000011010101001100000100",
"00111110000001000000000000100100",
"01010011000011010000011010110110",
"01010011000001000000000000100100",
"00000000001001001001000100001101",
"00000110101010000011111000000100",
"00000000001001001001010100001101",
"10100111000011010101001100000100",
"00111110000001000000000000100100",
"10100000000011010000011010011010",
"01010011000001000000000000100100",
"00000000001001001011001000001101",
"00000110100011000011111000000100",
"00000000001001001010110100001101",
"11001110000011010101001100000100",
"00111110000001000000000000100100",
"10110111000011010000011001111110",
"01010011000001000000000000100100",
"00000000001001001101100100001101",
"00000110011100000011111000000100",
"00000000001001001101001000001101",
"11100011000011010101001100000100",
"00111110000001000000000000100100",
"11011110000011010000011001100010",
"01010011000001000000000000100100",
"00000000001001001110110000001101",
"00000110010101000011111000000100",
"00000000001001001110011100001101",
"00001100000011010101001100000100",
"00111110000001000000000000100101",
"11101111000011010000011001000110",
"01010011000001000000000000100100",
"00000000001001010001011100001101",
"00000110001110000011111000000100",
"00000000001001010001000000001101",
"00100111000011010101001100000100",
"00111110000001000000000000100101",
"00011101000011010000011000101010",
"01010011000001000000000000100101",
"00000000001001010011011100001101",
"00000110000111000011111000000100",
"00000000001001110001010100001101",
"11011001000011010101001100000100",
"00111110000001000000000000100111",
"01111111000011010000011000001110",
"01010011000001000000000000100111",
"00000000001010000000110000001101",
"00000110000000000011111000000100",
"00000000001010000001010000001101",
"10110000000011010101001100000100",
"00111110000001000000000000101000",
"01001000000011010000010111110010",
"01010011000001000000000000101000",
"00000000001010001110011100001101",
"00000101111001000011111000000100",
"00000000001010001011011000001101",
"11111011000011010101001100000100",
"00111110000001000000000000101000",
"11101100000011010000010111010110",
"01010011000001000000000000101000",
"00000000001010010001001100001101",
"00000101110010000011111000000100",
"00000000001010010000000100001101",
"00101100000011010101001100000100",
"00111110000001000000000000101001",
"00011010000011010000010110111010",
"01010011000001000000000000101001",
"00000000001010010100001100001101",
"00000101101011000011111000000100",
"00000000001010010011101100001101",
"01010110000011010101001100000100",
"00111110000001000000000000101001",
"01001111000011010000010110011110",
"01010011000001000000000000101001",
"00000000001010011000000100001101",
"00000101100100000011111000000100",
"00000000001010010101110100001101",
"10010011000011010101001100000100",
"00111110000001000000000000101001",
"10001001000011010000010110000010",
"01010011000001000000000000101001",
"00000000001010011111000100001101",
"00000101011101000011111000000100",
"00000000001011011101111100001101",
"11100100000011010101001100000100",
"00111110000001000000000000101101",
"11100001000011010000010101100110",
"01010011000001000000000000101101",
"00000000001011011110101100001101",
"00000101010110000011111000000100",
"00000000001011011110100100001101",
"11110010000011010101001100000100",
"00111110000001000000000000101101",
"11110000000011010000010101001010",
"01010011000001000000000000101101",
"00000000001011011111100100001101",
"00000101001111000011111000000100",
"00000000001011011111011100001101",
"00111011000011010101001100000100",
"00111110000001000000000000101110",
"01100110000011010000010100101110",
"01010011000001000000000000101110",
"00000000001011101101111100001101",
"00000101001000000011111000000100",
"00000000001011101110101100001101",
"11111001000011010101001100000100",
"00111110000001000000000000101110",
"11110100000011010000010100010010",
"01010011000001000000000000101110",
"00000000001011110010100000001101",
"00000101000001000011111000000100",
"00000000001011110000011000001101",
"01111011000011010101001100000100",
"00111110000001000000000000101111",
"00110011000011010000010011110110",
"01010011000001000000000000101111",
"00000000001011111101000000001101",
"00000100111010000011111000000100",
"00000000001011111000100000001101",
"11100001000011010101001100000100",
"00111110000001000000000000101111",
"11011111000011010000010011011010",
"01010011000001000000000000101111",
"00000000001100000000111000001101",
"00000100110011000011111000000100",
"00000000001011111110110000001101",
"00111000000011010101001100000100",
"00111110000001000000000000110000",
"01000010000011010000010010111110",
"01010011000001000000000000110000",
"00000000001100001000001000001101",
"00000100101100000011111000000100",
"00000000001100000100110000001101",
"11011010000011010101001100000100",
"00111110000001000000000000110000",
"11100101000011010000010010100010",
"01010011000001000000000000110000",
"00000000001100010100001000001101",
"00000100100101000011111000000100",
"00000000001100010101010000001101",
"10011110000011010101001100000100",
"00111110000001000000000000110001",
"01111001000011010000010010000110",
"01010011000001000000000000110001",
"00000000001100011101011000001101",
"00000100011110000011111000000100",
"00000000001100011010111100001101",
"00000010000011010101001100000100",
"00111110000001000000000000110010",
"11100011000011010000010001101010",
"01010011000001000000000000110001",
"00000000001100100011011100001101",
"00000100010111000011111000000100",
"00000000001100100001000000001101",
"10000110000011010101001100000100",
"00111110000001000000000000110010",
"01000011000011010000010001001110",
"01010011000001000000000000110010",
"00000000001100101101101100001101",
"00000100010000000011111000000100",
"00000000001100101001001000001101"
)
,(
"11101011000011010101001100000100",
"00111110000001000000000000110010",
"11101000000011010000010000110010",
"01010011000001000000000000110010",
"00000000001100110011100000001101",
"00000100001001000011111000000100",
"00000000001100101111100100001101",
"10000000000011010101001100000100",
"00111110000001000000000000110011",
"10001101000011010000010000010110",
"01010011000001000000000000110011",
"00000000001100111001101100001101",
"00000100000010000011111000000100",
"00000000001100111001010000001101",
"00000011000011010101001100000100",
"00111110000001000000000000110100",
"10101010000011010000001111111010",
"01010011000001000000000000110011",
"00000000001101000010110100001101",
"00000011111011000011111000000100",
"00000000001101000001000100001101",
"01011111000011010101001100000100",
"00111110000001000000000000110100",
"00111101000011010000001111011110",
"01010011000001000000000000110100",
"00000000001101001000011000001101",
"00000011110100000011111000000100",
"00000000001101000110010100001101",
"10111011000011010101001100000100",
"00111110000001000000000000110100",
"10001101000011010000001111000010",
"01010011000001000000000000110100",
"00000000001101001111010000001101",
"00000011101101000011111000000100",
"00000000001101001100101000001101",
"00110001000011010101001100000100",
"00111110000001000000000000110101",
"01100000000011010000001110100110",
"01010011000001000000000000110101",
"00000000001101110100010000001101",
"00000011100110000011111000000100",
"00000000001101011110101100001101",
"10110000000011010101001100000100",
"00111110000001000000000000110111",
"01010001000011010000001110001010",
"01010011000001000000000000110111",
"00000000001101111110100100001101",
"00000011011111000011111000000100",
"00000000001101111100000000001101",
"00011110000011010101001100000100",
"00111110000001000000000000111000",
"11110100000011010000001101101110",
"01010011000001000000000000110111",
"00000000001110011110011000001101",
"00000011011000000011111000000100",
"00000000001110011110101000001101",
"00011100000011010101001100000100",
"00111110000001000000000000111010",
"00100110000011010000001101010010",
"01010011000001000000000000111010",
"00000000001110101000011000001101",
"00000011010001000011111000000100",
"00000000001111001101101000001101",
"00011001000011010101001100000100",
"00111110000001000000000000111101",
"00001100000011010000001100110110",
"01010011000001000000000000111101",
"00000000001111010111111000001101",
"00000011001010000011111000000100",
"00000000001111010010100000001101",
"10100110000011010101001100000100",
"00111110000001000000000000111101",
"10001000000011010000001100011010",
"01010011000001000000000000111101",
"00000000001111011101011100001101",
"00000011000011000011111000000100",
"00000000001111100000100000001101",
"00100100000011010101001100000100",
"00111110000001000000000000111111",
"10001010000011010000001011111110",
"01010011000001000000000000111110",
"00000000001111110101000000001101",
"00000010111100000011111000000100",
"00000000001111110010101000001101",
"01101110000011010101001100000100",
"00111110000001000000000000111111",
"01011000000011010000001011100010",
"01010011000001000000000000111111",
"00000000001111111001111100001101",
"00000010110101000011111000000100",
"00000000001111110111111000001101",
"10111011000011010101001100000100",
"00111110000001000000000000111111",
"10101101000011010000001011000110",
"01010011000001000000000000111111",
"00000000001111111101101000001101",
"00000010101110000011111000000100",
"00000000001111111100100100001101",
"11110000000011010101001100000100",
"00111110000001000000000000111111",
"11100010000011010000001010101010",
"01010011000001000000000000111111",
"00000000010000000010100000001101",
"00000010100111000011111000000100",
"00000000010000000010111100001101",
"00110100000011010101001100000100",
"00111110000001000000000001000000",
"00110001000011010000001010001110",
"01010011000001000000000001000000",
"00000000010000000100100000001101",
"00000010100000000011111000000100",
"00000000010000000100011000001101",
"01011101000011010101001100000100",
"00111110000001000000000001000000",
"01011011000011010000001001110010",
"01010011000001000000000001000000",
"00000000010000001000001100001101",
"00000010011001000011111000000100",
"00000000010000000110110000001101",
"10011111000011010101001100000100",
"00111110000001000000000001000000",
"10010001000011010000001001010110",
"01010011000001000000000001000000",
"00000000010000001011110000001101",
"00000010010010000011111000000100",
"00000000010000001011010000001101",
"00011000000011010101001100000100",
"00111110000001000000000001000001",
"01000000010001100000001000111010",
"01001111000011010101010100001000",
"00111110000001000000000001000001",
"10001100010001100000001000101110",
"01001010000011010101010101011010",
"00111110000001000000000001000001",
"01000000010001100000001000100010",
"01000101000011010101010100001001",
"00111110000001000000000001000001",
"01001000010001100000001000010110",
"01000000000011010101010100001001",
"00111110000001000000000001000001",
"01001100010001100000001000001010",
"00111010000011010101010100001001",
"00111110000001000000000001000001",
"01010101010101100000000111111110",
"00000000010000010010111100001101",
"00000001111101000011111000000100",
"00001101010101010000001001011010",
"00000100000000000100000100100101",
"01000110000000011110100100111110",
"00001000000000101111111111010100",
"00000000000000000000110101010110",
"00010100000000000000100000000000",
"01000110001011111101111100111110",
"00001000000000101111111111010100",
"11110000000000001000110111010110",
"10010100100000000000011111111111",
"01000110000001000100000001000110",
"01000110000000010000100101000000",
"01000100010001100000010000000000",
"01000110010101100000000100001001",
"01010101000000010000101001001100",
"00000001000010100101000001000110",
"00001001010010000100011001010110",
"01001100010001100101011000000001",
"01000110010101100000000100001001",
"01000110000000010000101001010100",
"01000100010001100000010000000000",
"01000000010001100000000100001001",
"00001001010000000100011000000100",
"00000000000100000100011000000001",
"00001001100100001001000101010110",
"11111111110110000100011000001110",
"10111000101011011001100000000001",
"11111111111101001100001010011111",
"00001010100000000100011010001001",
"01010110000001000000000001000110",
"01000000000010011001000010010001",
"00001111010101100000000000000101",
"10101101100110000001110100000001",
"11110101110000101001111110111000",
"00001101000010001000100111111111",
"00000100000000000010010100111110",
"00000011010001000011111001001000",
"00000000001001010010110000001101",
"00111011001111100100011100000100",
"01000000110010000000110100000011",
"00111110010010010000010000000000",
"10000000000011010000001100110010",
"01010110000001000000000000001110",
"01000110000000110010100100111110",
"01000110000000101111111111010000",
"01000110000111000001111111111110",
"00111110000000011111111111010000",
"01000110010101100001111000110101",
"01010101000000010000101001001000",
"00000001111111111101010001000110",
"00001000000111010000000100111110",
"00000010111111111110110001000110",
"00000001010110100001101000011010",
"00000000000011100001001000001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"01000110000001001000111100111110",
"00001000000000101111111111010100",
"00000010000010100100100001000110",
"00001110000101110000111000001110",
"00000001000010100100100001000110",
"11111111110101000100011000011000",
"11111111010001100000000000000001",
"00001010001011000010110100000000",
"00001000000000000000011101000010",
"01000000111101001110000100111110",
"01000110000000000000000011011100",
"00101100001011010000000011111110",
"00000000000011000100001000001010",
"01111000010001100101011000001000",
"00001110001111100000000100001010",
"00000000110001100100000000100001",
"00000000111111010100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"10110101010000000010100000110000",
"11111100010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000100001000010",
"00001000000111001000100100111110",
"00000000000000001010001101000000",
"00101101000000001111101101000110",
"00000111010000100000101000101100",
"10101001001111100000100000000000",
"00000000100100100100000000000010",
"00000000111110100100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"10000001010000000001110000110011",
"11111001010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000011101000010",
"01000000001101000011100000111110",
"01000110000000000000000001110000",
"00101100001011010000000011111000",
"00000000000001110100001000001010",
"00101110010000100011111000001000",
"00000000000000000101111101000000",
"00101101000000001111011101000110",
"00000111010000100000101000101100",
"01000101001111100000100000000000",
"00000000010011100100000000101110",
"00000000111101100100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"00111101010000000010111001010000",
"11110101010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000011101000010",
"01000000000000011100101100111110",
"01000110000000000000000000101100",
"00101100001011010000000011110100",
"00000000000001110100001000001010",
"00100001000110010011111000001000",
"00000000000000000001101101000000",
"00101101000000001111001101000110",
"00010000010000100000101000101100",
"00000000000011010000100000000000",
"01000110100000000000000000000000",
"00111110000000010000101001111000",
"00000001010000000010000001001001",
"11101100010001100000100000000000",
"00000001010110100000001011111111",
"00111101111111101111010001000000",
"11111111111111111101100010001101",
"11010011100000101000111000000101",
"10001110100101111001101010011010",
"00010000100111010000000100010000",
"10001000000100001001110100000001",
"10001000100000011000111100000001",
"01001101000000000000110000111101",
"01001001010011000100110001001001",
"01001111010000110100010101010011",
"00001001010100110100010001001110",
"01000101010100100101000000000000",
"01001001010100110100100101000011",
"00000000000010010100111001001111",
"01010101010001000100111101001101",
"01001111010101000100010101001100",
"01000100000000000000011101010000",
"01010100010101000100001101001001",
"00000000000001000101000001001111",
"01000101010100110100000101000010",
"01010000010100110000000000000100",
"00000000000001000100111001000001",
"01000101010100100100010101001000",
"00011001000011100001111000001110",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"10010001010101100001111000001010",
"00000100000011110000100110010000",
"00110101000101110000010000001111",
"00001010000000000000010001000010",
"00001000001111011000100100001010",
"00011000000010001001000000011000",
"10101101100110001000100000010000",
"11100101110000101001111110111000",
"01010110000010011000100111111111",
"01100011000000000000011000111101",
"01110100011000010110010101110010",
"00000000000000000000110101100101",
"11011000000011010000011000000000",
"00000010000001011111111111111111",
"01000000000010011001000010010001",
"00010001100100000000000000101000",
"11111111010001100000001000011101",
"00101101000100000001110000000000",
"10001000000100000000101000101100",
"01000010000111000010001000101100",
"00010000000011110000000000001110",
"11111111100111000011111000000010",
"00000000000001000100001000101100",
"00111101100010010001000000001001",
"10010000000110100001101001010011",
"10111000101011011001011000001000",
"11111111110100101100001010011111",
"00010111000011100000100010001001",
"00111110010101100000111000111101",
"01000010001101011111111110110111",
"00110101000010100000000000000010",
"11111111111100010011111000111101",
"01010110000000000000010001000010",
"00001000000000010001110100001111",
"00000000000000000000010000001101",
"00000000000000000000110100000110",
"11011000000011010000011000000000",
"00000010000001011111111111111111",
"00001001100100001001000100011101",
"00010000000000000001000101000000",
"00000000000001100100001000000010",
"01000000100010010001000000001000",
"00011010010100110000000000001101",
"10010110000010001001000000011010",
"11000010100111111011100010101101",
"01010101100010011111111111101001",
"00001101000101110001101000011010",
"00000101111111111111111111011000",
"00000000000001000011110100000001",
"01000100010011100100100101000110",
"10010000000111010000111100110110",
"00000000111111110100011000000010",
"10000010100111010001110000011100",
"00101100001011010101011000000000",
"00000000000001110100001000001010",
"00111101100010000000100000001000",
"00000000000000000011111101000000",
"00001010001011000010110101010011",
"00001000000000000000011001000010",
"00110001010000000011110100001000",
"00101101010100010000000000000000",
"00010100010000100000101000101100",
"11001100100011010000100000000000",
"10000001000001011111111111111111",
"00001101000111010001110100011101",
"00000101111111111111111111011000",
"00010101010000000011110100000001",
"00101101010100000000000000000000",
"00001100010000100000101000101100",
"11111100100011010000100000000000",
"10000001000001011111111111111111",
"00000001010000000011110100001000",
"00010000000010000000100000000000",
"00000000000001100011110110001000",
"01100111011100100110111101100110",
"00111110010101110111010001100101",
"00101100000010100010001010110111",
"00000000000010110100001010010000",
"11110000001111100101000100001110",
"10011100100100000011010111111110",
"00001000111111111000010100111110",
"11000010000000100010110000111110",
"00010010000011010000000000001000",
"01000000000001000000000000001110",
"00001001000011010000000000000101",
"00111110000001000000000000001110",
"00001110000111100000001000011001",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000001101101100011111000100010",
"01000110000000000000011100111101",
"01000101010011000100100101000001",
"00000000000000110011111001000100",
"00000111001111100100101101001111",
"01000101010110000100010100000000",
"01000101010101000101010101000011",
"00011010000110100001110001000111",
"00011100010001110011110100000001",
"00111101000000100001101000011010",
"01000101010100110000000000001001",
"01000011010001010101011001010100",
"00111110010100100100111101010100",
"00001001001111011111110000101001",
"01010100010001010100011100000000",
"01010100010000110100010101010110",
"01001111010001100101001001001111",
"00011110010000100000010000001010",
"00000011001111100100011100000000",
"00000000000101000100011000000001",
"01010110000000010011100100111110",
"01000110001000101101000100111110",
"11110011001111100000000000011001",
"00001010011011000100011000000000",
"11111111111111000000110100000010",
"00111110000000010000010111111111",
"00000100001111011111101111100101",
"01001001010101010101000100000000",
"00000001000011100101101001010100",
"01000001000000000000010100111101",
"01010100010100100100111101000010",
"00000010111111111101010001000110",
"00000000000011101100101100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00001101000000010010011100111110",
"00000101111111111111111111100100",
"00000000000100000100011000000010",
"11111111111111111110010000001101",
"00111110000100000000000100000101",
"11100100000011010001011000000011",
"00000001000001011111111111111111",
"11111111110110000100011000001110",
"11111111110101000100011000000001",
"01000010010000000000110100000001",
"10010001010101100000000000001111",
"10101101100110000000100110010000",
"11111001110000101001111110111000",
"00100011001111011000100111111111",
"01100100011011100111010100000000",
"01101110011010010110011001100101",
"01101001001000000110010001100101",
"01110010011101000111001101101110",
"01101001011101000110001101110101",
"01101100001000000110111001101111",
"01110100011000010110001101101111",
"01101110001000000110010001100101",
"00100000011100100110000101100101",
"01001111010100110000000000000111",
"01001110010010010101010001000110",
"11111111110101001100011001010100",
"00001010010001001100011010000010",
"00011000010001101000001010001110",
"11111111111011000100011000000000",
"00010111000111000000111100000010",
"00011100001101100001000000101100",
"10011001000000000010101001000010",
"00001010010000000100011010011001",
"01000110000111100000111000000010",
"01000110000111000000001111111111",
"01000110000000010000101001000000",
"00001110000101100000000001000000",
"00000100000110000000111100000100",
"00001010001000100010000001001110",
"00000001111111111110000001000110",
"00000010111111111110110001000110",
"11000101010000000000000101011010",
"10001000100000011000111111111111",
"10000001111111111101010011000110",
"01011010000000001000000001000110",
"01000100010001100011110100000001",
"00000000010001100000001000001010",
"00111101001010100001011100000100",
"01000010111111111111001100111110",
"11010100110001101111111111111010",
"01000100110001101000001011111111",
"01000110100000101000111000001010",
"00010000000000100000101001000000",
"00000011111111110100011000010110",
"00000000010000000100011000011100",
"00100011010011100000111100010110",
"00000011000000110001100000001111",
"10001000100000011000111110011110",
"10000001111111111101010011000110",
"01000110111111110111011000111110",
"00000001010110100000000001000000",
"01000101000000000000010100111101",
"00111111010101000100100101001101",
"00011100000000001111111101000110",
"00000000000110110100011000001110",
"01000010000111110011100000010111",
"00000000010001100000000000000100",
"10101111001111100010001000000001",
"10010001010101100011110111111111",
"00000111010000000000100110010000",
"00111110000001000000111000000000",
"10011000000110001111111111011110",
"11000010100111111011100010101101",
"00001000100010011111111111110011",
"00111110010101100011110100000001",
"11100001001111101111111110010010",
"00000000000110100100011011111111",
"00111101111111111000100100111110",
"11111111100001000011111001010110",
"01000110111111111011110100111110",
"01111011001111100000000000011010",
"00000000000001000011110111111111",
"01000101010100000101100101010100",
"11111111011100000011111001010110",
"00001001100100001001000101010110",
"01000110000000000000011101000000",
"10011111001111100000000000100000",
"10111000101011011001100011111111",
"11111111111100111100001010011111",
"00000000000110100100011010001001",
"00111101111111110101010100111110"
)
,(
"01001101010001010000000000000100",
"00111110010101010101010001001001",
"00000110001111011111111111010110",
"01000001010100000101001100000000",
"01010110010100110100010101000011",
"01001001111111110011110100111110",
"01001100111111110111010100111110",
"01000110111111110111000100111110",
"00101111001111100000000000011010",
"00000000000001010011110111111111",
"01000011010000010101000001010011",
"00110100001111100101011001000101",
"11111111100010100011111000100100",
"00100100001011010011111001010111",
"01000011000000000000001000111101",
"00100010000011110000111101010010",
"00000000000010000100001000101100",
"00001110000010100000101000001000",
"00111101000011100001100100001110",
"10010000100100011001100011010110",
"00010001000011110000111100001001",
"00010111000010101001000100010000",
"00100110000010101001000100010000",
"00010001000010011000100100010000",
"00010001000111110100001100010000",
"00011100000111110010101010001001",
"10010000000000000000101001000010",
"00100101000011101001101000001000",
"11011000010000001000100000010000",
"11010110100010000001000011111111",
"00100110010000100011010110001110",
"00001000100100000001100100000000",
"00001010100100011001000010010001",
"00001010100100010001000000010111",
"01000011100010010001000000100110",
"00000000001101100100001000011111",
"00010000001000110101010100010001",
"00010000100010010010100001010101",
"10001110000110101000100100010001",
"00001000100100000001100010100101",
"00001000111111111101011001000000",
"00000000001101100100000000001001",
"00000000001010000100001000110101",
"00001001100100011001000000011001",
"10001000000100000010001101010101",
"10010000100100010010100001010101",
"00010000000101100000101010010001",
"00010000001001010000101010010001",
"01000010000111110100001110001001",
"00010000000100011111111111001010",
"10001001000100010001000010001001",
"10010000101001011000111000011010",
"11111111110101000100000000001000",
"00010110000010101001000100001000",
"00100101000010101001000100010000",
"00010000000100011000100100010000",
"00000000000001010011110110001001",
"01001110010010010101001001010000",
"00010111000011101001000001010100",
"01001100001111101000100000010000",
"00001001100100001001000111111111",
"10001001000100000001000100001010",
"01010101000000000000011100111101",
"01001101010001000010111101000100",
"11100100001111100100010001001111",
"00000110001111010000101011111111",
"00101111010001000101010100000000",
"10010000010001000100111101001101",
"00101010000011111001000100001000",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00000001010000100010100100010001",
"11011001001111100010000100000000",
"11000010101010101010010011111111",
"10010000001000010000000000000110",
"10001000000100000010000100001000",
"01010101000000000000011000111101",
"01001111010011010010111101001101",
"11001110001111101001000001000100",
"00101001000010001001000011111111",
"00010001000000000000100101000010",
"00000000000000010100001000101010",
"10011001000101100001000100100001",
"00000110001111011000100100010000",
"00101111010011010101001100000000",
"10010001010011010100010101010010",
"00010000010101100000100110010000",
"00000000000000010100001000101001",
"01000010001010010001000100100001",
"10100100001000010000000000000001",
"01010110000000000010000001000110",
"10010001000010011001000010010001",
"00100110000011100001101110010000",
"00101000010101010001011000011100",
"00101000010101010001000000010001",
"10111000101011011001100010001001",
"11111111111010111100001010011111",
"11000010101010100000101010001001",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"00111101100010000001000000001010",
"01001101010001100000000000000110",
"01000100010011110100110100101111",
"00001010111111111011100000111110",
"01001101000000000000001000111101",
"10010000000010001001000000101010",
"00010000100010000001000000101010",
"11111111010110110011111010001000",
"00101010000000000000000100111101",
"00001010111111111110111000111110",
"00101111000000000000010000111101",
"00111110010001000100111101001101",
"00111101000010001111111111100011",
"10010000001011110000000000000001",
"11111111100010110011111000001000",
"00111010001111101000100000010000",
"00000000000000110011110111111111",
"00111110010001000100111101001101",
"00111101000010101111111111101101",
"00101111001010100000000000000101",
"00001111010001000100111101001101",
"00000000001011010100011000000100",
"01000010000010100010110000101101",
"10001110110101110000000000000101",
"11010110000000000000011101000000",
"00000000001010111100011010010000",
"11000010000010001010110010010111",
"10010000000110010000000000000110",
"10001000000100000001100000001000",
"11000010101101110000100010010000",
"00000100100100000000000010010011",
"00101101000000000011000001000110",
"01000110000011110000101000101010",
"00111000000101110000000000111001",
"00110000010001100001111100100010",
"01000110000101110001110000000000",
"00101010001011010000000001000001",
"01011010010001100000111100001010",
"00100010001110000001011100000000",
"00000000001101110100011000011111",
"01100001010001100001011100011100",
"00001010001010100010110100000000",
"00000000011110100100011000001111",
"00011111001000100011100000010111",
"00011100000000000101011101000110",
"11111111111001000000110100010111",
"00101101000000100000010111111111",
"00000110010000100001111100101010",
"10001000000100000000100100000000",
"10010001000000000100011001000000",
"10010000100100010000100110010000",
"00010001000011100101011000001001",
"11000010101101011000100100010000",
"00001110100110110000000000100011",
"00001110010000100010011000001110",
"10010001100100001001000100000000",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00001111100010010001000000010001",
"00010110000010101001000100001111",
"00100101000010101001000100010000",
"11011001010000001000100100010000",
"00010001000100000000100111111111",
"00010110000010101001000110001001",
"00100101000010101001000100010000",
"10001000000100001000100100010000",
"01101001010000001001100100011000",
"10010001100010100001000111111111",
"00000000000010010100001000001010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"10001001000100010001000010001000",
"00101010000000000000001000111101",
"00011001000011100001111000101111",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00001000111111110010000000111110",
"00111110000000000000011100111101",
"01000010010011010101010101001110",
"01000010001010010101001001000101",
"00111110001000010000000000000111",
"01000111010000000000000001010100",
"00000000010000000100011000000000",
"00000100010000100011100000101101",
"00010000000010101001000100000000",
"00001000100100000000100010001000",
"10001010000100011010101010010001",
"00101101000000000001111101000110",
"00000000000011100100001000111000",
"00001001100100000001100100010111",
"00010000000010101001000100010001",
"01000000100010000001000010001000",
"10010000000010001111111111101010",
"00100000010001100000111100100011",
"00100000000101110001000000000000",
"00010000000010101001000100100010",
"00010001001000110001000010001000",
"00010000000000000010000001000110",
"00100010001000000001011110001001",
"10001000000100000000101010010001",
"01000011000000000000011100111101",
"01000101010101100100111001001111",
"01000010001010010101010001010010",
"00111110001000010000000000000111",
"00111011010000001111111110011100",
"00000000010000000100011000000000",
"00000100010000100011100000101101",
"00010000000010101001000100000000",
"00011111010001100000100010001000",
"01000010001110000010110100000000",
"00011001000101110000000000001111",
"00001010100100010000100010010000",
"00010111000011101000100000010000",
"11101001010000001000100000010000",
"10010001100100000000100011111111",
"00010000000010101001000100100000",
"00010000001000000001000110001000",
"00010001000000000010000001000110",
"10010001001000100010001100010111",
"10001001100010000001000000001010",
"01000001000000000000011000111101",
"01000110010010010100100001010011",
"00000111010000100010100101010100",
"10101001001111100010000100000000",
"00000000001110100100000011111111",
"00101101000000000100000001000110",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"00000000000111110100011000001000",
"00001111010000100011100000101101",
"10010000000110010001011100000000",
"10010001000101110000111000001000",
"00010000100010000001000000001010",
"11111111111010010100000010001000",
"00001111001000111001000000001000",
"00010000000000000010000001000110",
"10010001001000100010000000010111",
"00010000100010000001000000001010",
"00001010100100010010001110001000",
"00000110001111011000100000010000",
"01001001010010000101001100000000",
"10010001010011000101010001000110",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10010000100100011000100000010000",
"00101010000011111001000100001001",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"10001010000100011000101000010001",
"10010000000010011001000110010000",
"00001110010101100000100110010001",
"00110101000000000100000001000110",
"00011001000000000011010001000010",
"10010000000110100000100010010000",
"00010000001001010000111000001000",
"00010001100010100001000110001000",
"00010000100110101000100100010000",
"10010000101001011000111010001000",
"00001000100100001001000100001000",
"10010000100010100001000110010001",
"00001100010000100100001100001000",
"00010110000010101001000100000000",
"00100101000010101001000100010000",
"00000001010000001000100100010000",
"10001000000100000000100100000000",
"00001000111111111100100001000000",
"10101010101001001000100110001001",
"00100001000000000000100111000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"01010011000000000000011000111101",
"01010100010001100100100101001000",
"00101010000011111001000101010010",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"10010001000010011001000110010000",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10001010000100011000100000010000",
"00111110101001001000101000010001",
"11000010101010101111101111000111",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"10010000100010000001000000001010",
"00010000000010100000101000001000",
"00000000000000100011110110001000",
"00001111100100010010101001000100",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00001001100100011001000010001000",
"01000010001010100000111110010001",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"00010001100010000001000000001010",
"10100100100010100001000110001010",
"00001001111110111000011000111110",
"00000000000010011100001010101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00000000000000100011110110001000",
"00001000100100000010111101000100",
"00000000000000000000000000001101",
"10001000000100000010010010000000",
"01000100000000000000010000111101",
"00001111010001000100111101001101",
"01000010001011000010001000001111",
"00001111001111010000000000000001",
"00000000000011110100001000101010",
"00100001000011000011111111000110",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"11000110000000000000001101000000",
"00001111100110010000010000111111",
"00010110000010101001000100001111",
"00100101000010101001000100010000",
"01000010010000111000100100010000",
"00100011010010101111111111110000",
"00000000000101000100011000001111",
"00001000100100000010001000100000",
"01000110000100010010001101001010",
"00100010001000000000000000010100",
"00000111001111011000100100010000",
"01000101010011100100011000000000",
"01000101010101000100000101000111",
"10010000100100010000100010010000",
"00000000000000000000110100001001",
"11010100010101100011111111110000",
"00101001100010000001000010001011",
"00100001000000000000000101000010",
"00000000001000100100001000001110",
"00001001010000100100001100011011",
"00001010100100010001000100000000",
"00000001000001110011111000010001",
"10001010000100011000100000010000",
"10001010000100010000101010010001",
"11111010001111100000111100001111",
"00010001000010101001000100000000",
"01000000000010101001000110001010",
"10001001000010001111111111011010",
"00000000000011111100001010101010",
"00001101000010011001000010010001",
"00111111111100000000000000000000",
"10001001000100000001000101010110",
"00111101000000110001011100111110",
"00111110010001000000000000000011",
"00001001100100011001000001000110",
"00010001000100000000111001010110",
"11111100010111110011111010001001",
"01000110000001000000111110010000",
"00101100000101110000000000101110",
"01000010000111000011011000001111",
"00011001100010000000000000110010",
"10010000000110000000100010010000",
"00101010000011111001000100001000",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00111110000100011000101000010001",
"00001000100100001111110000110101",
"00001010100100011000101000010001",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"10001001000100010001000010001000",
"10010000101000011001011110010000",
"00001010001111100000100110010001",
"01000110000001000001000011111111",
"00101100001011010000000001000101",
"01100101010001100000111100001010",
"00100010001011000001011100000000",
"00011100001101100001000100001010",
"01010110000000000001000001000010",
"00010001000110000001000000001110",
"11110110001111101000100100011001",
"10010110100100000000100111111011",
"10001001000010011001000110010000",
"11111111111001000000110101010110",
"00111110000000100000010111111111",
"10001000000100001111111011011001",
"00111110111111110010000100111110",
"00111101010101110000000001001001",
"01010110000000000011010101000110",
"10010001000010011001000010010001",
"10101000110101011001000010011011",
"00001001100100011001000000001001",
"00011011000010001001000011000011",
"00101000010101011000100000010000",
"00010001000000000000100011000010",
"00010001000010001001000000010110",
"00010000100010000001000000100101",
"00010000000100011000100100010001",
"10111000101011011001100010001001",
"11111111110101111100001010011111",
"10010000000010010000100110001001",
"10101000110101010001101100001000",
"00100101010101101010010111010110",
"00000110001111011000100000010000",
"01001100010001100011111000000000",
"10010000010101000100000101001111",
"11111111100011011001000000001000",
"10011100000000000000111111111111",
"11110000000000000000000000001101",
"00001101000011100001110011111111",
"01111111111100000000000000000000",
"00000110010000100011011000011100",
"00000000000000001000110100000000",
"10010001101000100000000000010000",
"00010000000010101001000100001010",
"00001111111111111111111110001101",
"00000000000011011001110000000000",
"00011100111111111111000000000000",
"00000000000000000000110100001110",
"00110110000111000111111111110000",
"10001101000000000000011001000010",
"00000000000100000000000000000000",
"10100100100100011001000010100010",
"00000000000000000000000010001101",
"00000000000011011001110010000000",
"00011100011111111111000000000000",
"00010000000010101001000100011011",
"00000000000000000000110110001000",
"00011011000111000111111111110000",
"00000000000000000000110100010110",
"00001101000101110001111111111000",
"00111111111100000000000000000000",
"01000010000010100011100000101101",
"10011010000010000000000000001110",
"11100000000000000000000000001101",
"01010110001010000101010111111111",
"00111101100010011000100110001000",
"00000000000001110100001000101001",
"10001000010101100001000000001000",
"00011010001111011000100110001001",
"01010110101000100000100010010000",
"00010001100010100001000100001110",
"10010001000011110000111110001010",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"10001010000100011000101000010001",
"00001111111111110001010100111110",
"00010000000000000000000000001101",
"00001010001010100010110100000000",
"10001101000000000000011001000010",
"10000000000000000000000000000000",
"11111111111111110000110110011100",
"00111000000101110000000000011111",
"10010000000000000000110101000010",
"10101000110101010001101100001000",
"00000000100011011000100000010000",
"10010110000000000001000000000000",
"11111111000011010000100010010000",
"00011100000000000000111111111111",
"10001001000100000010001000010001",
"00001000100100001001000100111101",
"00001111111111111111111100001101",
"00001101000100010001110000000000",
"01111111111100000000000000000000",
"00000110010000101001000000011100",
"00000000000000000000110100000000",
"00010001001000100000000000010000",
"00001000100100000001101010001010",
"10001000000100000010010100001110",
"00001001010000100010101000010001",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10001001000100001000100000010000",
"01000110000000000000001000111101",
"00000000001100100100011000101010",
"00001000100100000010101000010111",
"00010000000100010000101010010001",
"00010101010001100001101010001001",
"00001000100100000010001100000000",
"00010000000100010000101010010001",
"00010101010001100001101010001001",
"00001111000011110010001100000000",
"00000001010000100010100100010111",
"00110110010001100010000100000000",
"00001111001010100001011100000000",
"00001010000010100001110000110110",
"10010000100100010011110100011100",
"11111111100100010011111000001001",
"00001010100100011000101000010001",
"10001000001111101000101000010001",
"00010001000010001001000011111111",
"00100011000000000001010001000110",
"00000000000101000100011000010000",
"01000010001010010001011100100011",
"10010001100010100000000000001111",
"00100001000010101001000100001010",
"00010000111110110001001100111110",
"00000100010000001000100100010001",
"00001001001111101000100000000000",
"00010110000010101001000111111011",
"00100101000010101001000100010000",
"00001111100110101000100100010000",
"00001000101010001101010100011010",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"00001111000011111000100000010000",
"00000110010000100010110000100010",
"00000000000000001000110100000000",
"00001111100111001000000000000000",
"00100000000000000000000000001101",
"00010000001010100001011100000000",
"00010100010000100001110000011010"
)
,(
"10010001000011110000111100000000",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00010000000000000000000010001101",
"11011110010000001001011100000000",
"01010100100010000001000011111111",
"00001001100100001001000101010110",
"00001101000011110000100010010000",
"00000000001111111111111111111111",
"00011010000100000011100000010111",
"11100000000000000000000000001101",
"00011100001101100001011111111111",
"10010000000000000000110101000010",
"10001000000100000001101100001000",
"00000000100011010010100001010101",
"10010110000000000001000000000000",
"10010001000110000000111001010110",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"10001000000100000001110001011000",
"10011111101110001010110110011000",
"10001001111111111100010111000010",
"00001000100100000000100010010000",
"01010101100010000001000000011011",
"11111111000011010000111100101000",
"00010111000000000000111111111111",
"00101100000110100001000000111000",
"00000000000001100100001000011100",
"00010000000000000000000010001101",
"00001000100100001001011000000000",
"00001111111111111111111100001101",
"00100010000100010001110000000000",
"00111110001111011000100100010000",
"00001101001111101111110001000100",
"00000000000000100011110111111111",
"00011010000011110010101101000110",
"01000010001011000010001000001111",
"00001010000010000000000000001011",
"11111111111111110000110100100100",
"01010111001000100111111111111111",
"00001101000011100000111100111101",
"00000000000011111111111111111111",
"00000000000011010000111100011100",
"00011100011111111111000000000000",
"00001101000000000000011001000010",
"00000000000100000000000000000000",
"10010001100100000000101000100010",
"10010001000010001001000000001001",
"11111111100011011001000110010000",
"10011100000000000000111111111111",
"00000000000000001000110110010001",
"11000010100111000111111111110000",
"00000000100011010000000000000110",
"10100010000000000001000000000000",
"00010000000011100101011000001001",
"00011010000100001000100100010001",
"00100011000000000001010101000110",
"00010101010001100001101000010001",
"01000110000101110010001100000000",
"00001101000101100000001111111111",
"00000000000000010000000000000000",
"00000000100011011010010000010110",
"10011100100000000000000000000000",
"00001111101000100000100010010000",
"00010001100010000001000000001111",
"10010001000100010000101010010001",
"10010001000100000001011100001010",
"10001001000100000010011000001010",
"01000010000111110010101000001000",
"00010001000100000000000000001101",
"10100101100011100001101010001001",
"10011000000010011001000110010000",
"00010000111111111101110001000000",
"00000001111111111111111100001101",
"11111110000011010001110000000000",
"00101101000000000000000100000111",
"00001111010000100000101000111000",
"00001000000010010000100100000000",
"00000000000000000000110110011010",
"00101000010101011111111111100000",
"00111101100010001000100101010110",
"00000000111111111100101100001101",
"00001010001010100010110100000000",
"00001001000000000000111001000010",
"00000000100011010000100000001001",
"10011100100000000000000000000000",
"10001000100010010101011000010000",
"00000000000000000000110100111101",
"00101010001011010000000000000001",
"00000000000011010100001000001010",
"00000000000000000000000010001101",
"00000000010001101001110010000000",
"00000010010000000010001000000000",
"01000110000101110000111000000000",
"10001101000101100000000000110111",
"10000000000000000000011111111111",
"00010001100010000001000010011100",
"00010001000010101001000110001010",
"10010001000010001001000010001010",
"10110111100010100001000100001010",
"10011001000000000010100111000010",
"00001010100100011001000010010001",
"00001010100100010001000000010111",
"01000011100010010001000000100110",
"00000000001011010100001000011111",
"00001110000010001001000000011010",
"00011010000010001001000000100101",
"00100101000011100000100010010000",
"00010000100010000001100000010000",
"00010000000100011000100100010001",
"11111111110100110100000010001001",
"00000000001010001100001010110111",
"10010001100100001001000110011001",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"11010011010000100001111101000011",
"00001000100100000001101011111111",
"00001000100100000010010100001110",
"00001110000010001001000000011010",
"00010000100010000001000000100101",
"00010000000100011000100100010001",
"11111111110101000100000010001001",
"10010001000010010000100110001000",
"00011011000010001001000010010000",
"10100101110101101010100011010101",
"10001000000100000010010101010110",
"00000000000000000000110100001111",
"00001101000111000000000000110000",
"00000000000100000000000000000000",
"00000101010000100010110000010111",
"01000000100110011000100100000000",
"00010001000010010000000000001110",
"00100101010101101001011011010100",
"00011011101010001101010100011011",
"00101000010101011000100100010000",
"11111111000011010000100010010000",
"00011100000000000000111111111111",
"00000000000101010100011000010001",
"00001000000110100001000100100000",
"00010000001000100010100001010101",
"00000000000000100011110110001001",
"10010000100100010010110101000110",
"00001101000100010101011000001001",
"10000000000000000000000000000000",
"01000110000110100001000100011100",
"01000110001000110000000000010101",
"00011111000101110000001111111111",
"00010110000000111111111001000110",
"00100000000000000001010101000110",
"10010000001000100010001101010101",
"00010001000011110101011011010110",
"00000100001111100000101101010010",
"01000110000110100001000111111101",
"01000110001000110000000000010101",
"00101010000101110000011111111111",
"00000000001000100100001000011100",
"00111110100010010001000000010001",
"00001111000011111111110100100000",
"00001111000011110000111100001111",
"00010001111110111101010000111110",
"11111011110011110011111000010000",
"10010001111111011111110000111110",
"00001011010101000000100110010000",
"01000000000011000101010000011000",
"00001000100100001111111111001000",
"00010000000100010000101010010001",
"10001001100010010000100010001001",
"01000110000000000000001000111101",
"00000000000011010000111100101111",
"00011100100000000000000000000000",
"11100000000000000000000000001101",
"00111110010101100010001000111111",
"01111101001111101111110011100100",
"00000000000000000000000000000000",
"00000000000000000000110100001111",
"01000110000111000111111111110000",
"01000110001000110000000000010100",
"00101001000101110000001111111111",
"00001000000000000000011101000010",
"01000000000011100101011000001001",
"00111110010001100000000001010011",
"00001010001110000010110100000000",
"00001001000000000001011101000010",
"00000000000010010100001000101010",
"00000000000000000000000000001101",
"00000110010000000101011010000000",
"11111111111111110000110100000000",
"01000000010101110111111111111111",
"10010001100100000000000000110011",
"11111111000011011001000000001001",
"00011100000000000000111111111111",
"00010000000000000000000000001101",
"10001010000100010010001000000000",
"00000000001101000100011000010001",
"00000110010000100011011100010111",
"11111000000111100011111000000000",
"00100001000000000000010001000000",
"10101010111110000110011000111110",
"00100001000000000000100111000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00000000000010100011110110001000",
"01001001010000110100010101010010",
"01000011010011110101001001010000",
"00001101000011110100110001000001",
"01111111111100000000000000000000",
"00000000000000000000110100011100",
"00101001000101110011111111110000",
"00001001000000000000100101000010",
"00000000000000000000000000001101",
"00111101010101100001110010000000",
"00100011000000000001010001000110",
"10010000000000000011010011000110",
"11000010101101111001011100001000",
"11000110010101110000000000011000",
"10101001100101110000000000100000",
"01000110000000000000101011000010",
"00010110000100000000000000100000",
"00000101010000000001110000100000",
"00100000000100000000101000000000",
"00111101100010000101011000011100",
"00111110010001100000000000000011",
"00111110000011110000111101000100",
"10010000100100011111111110110100",
"00001010100100010000100010010000",
"10001000000100001010010000100100",
"00010001000111110010110000100010",
"10001010000100010001110000101010",
"10001010000100010000101010010001",
"00001101000000000000100111000010",
"00111111111100000000000000000000",
"11111100111000110011111001010110",
"01110011000000000000011000111101",
"01110000011010010111001001110100",
"01010001000011110000111101100110",
"00111110000010110101000100001011",
"00011010000011111111110011010001",
"00101010000011110011011000100010",
"01000010000111110000101000011100",
"10010000100100010000000000001001",
"00010000000100010000100100001001",
"00001001000011110000111110001001",
"01000110000000000000010100111101",
"01010010010011110100111101001100",
"00001011010100010000111100001111",
"10101010001111100000101101010001",
"00100010000110100000111111111100",
"00011100001010100000111100110110",
"00000000000010010100001000001010",
"00001001000010011001000010010001",
"00001111100010010001000000010001",
"00000100001111010000100100001111",
"01000001010011010100011000000000",
"00111110000011110000111101011000",
"10010000100100011111111100111000",
"00001010100100010000100010010000",
"10001000000100001010010000100100",
"00010001000111110010110000100010",
"00010001000111000001111100101010",
"00010001000010101001000110001010",
"00000000000010011100001010001010",
"11110000000000000000000000001101",
"01111001001111100101011000111111",
"00000000000001000011110111111011",
"01001110010010010100110101000110",
"00111110000010011001000010010001",
"00010000000100010000001000101110",
"11111010001000110011111010001001",
"00111101000000011100100000111110",
"01010010010001100000000000000110",
"01000100010011100101010101001111",
"00001101000000000101000000111110",
"00111111111110010010000111111011",
"01000100001011010001100000001101",
"11111100001101110011111001010100",
"00111101111110000111101100111110",
"00101010010001100000000000000011",
"00001111000011110000111100101010",
"11111001111101110011111000001111",
"11110000000000000000000000001101",
"00011110001111100101011000111111",
"00000011010001000011111011111100",
"00111110111110110010101100111110",
"00000101001111010000000111101010",
"01000011010000010100011000000000",
"10110001000011010101001101001111",
"00001101010000000000001001101011",
"10111011101101010101010100010111",
"00111110111110011101000000111110",
"00000110001111010000000101110101",
"01000011010000010100011000000000",
"10010001010010000101001101001111",
"00000000000000000000110110010000",
"00010001010101100011111111110000",
"00001111000011111000100100010000",
"00111110111110011011010000111110",
"00000111001111101111101111100001",
"11111011111001100011111000000011",
"00111101000000000010100100111110",
"01000001010001100000000000000101",
"00001111010001110100111101001100",
"00111110000011110000111100001111",
"00000000000011011111100110011001",
"01010110001111111111000000000000",
"00111110111110101101001100111110",
"11001101001111100000001011100110",
"00000001100011000011111011111010",
"01000110000000000000010100111101",
"01001110010010010101001101000001",
"00001111000011110000111100001111",
"00111110111110010111100000111110",
"10010000100100011111011111101100",
"00001001100100001001000100001001",
"00001111000100000001000101010110",
"00111110000010110101001000010001",
"00100010010000101111101001110111",
"10001001000100000001000100000000",
"01011010001111100001000000010001",
"01010010100100001001000111111001",
"01010001000011100001100000001011",
"10010000000110000001101000001100",
"00111110100010000001000000101010",
"10000001001111101111011111010001",
"11111010100001100011111011111011",
"10010000111111111101010001000000",
"00010001000010101001000100001000",
"10001001000010001000100100010000",
"00000000000001100011110110001001",
"01001001010100110100000101000110",
"00001011010100110100100001001110",
"00111110100100010000100010010000",
"10100011001111101111101101100000",
"00010111110000101010101011111111",
"00100001111110110000110100000000",
"00011000000011010100000000001001",
"10101001010101000100010000101101",
"00111110000000000000011011000010",
"00000011010000001111101100111101",
"11111010010010100011111000000000",
"00000000000001010011110110001000",
"01000001010101000100000101000110",
"00000000000000000000110101001110",
"00111110010101100011111111110000",
"00001111000011111111101000111000",
"00000000000000000000000000001101",
"00011010001111100101011001000000",
"11110111010111100011111011111011",
"00111110111110110001111100111110",
"00000000000011010000000011100110",
"01010110001111111110000000000000",
"00111101111110001101100000111110",
"01000001010001100000000000000110",
"00110010010011100100000101010100",
"11001010001111100000111100001111",
"11110111001111100011111011111000",
"01010110000010011001000010010001",
"11110000000000000000000000001101",
"10010000100100010101011000111111",
"00001011010100100001000100001111",
"01000010111110011100011000111110",
"00010000000100010000000000100010",
"00111110000100000001000110001001",
"00001011010100101111100010101001",
"00001100010100010000111000011000",
"00111110000110010000111000011010",
"00100010001111101111001110100101",
"11111010110100100011111011110111",
"11010101001111101001000010010001",
"11111111110101000100000011111001",
"00001010100100010000100010010000",
"00001000100010010001000000010001",
"00000110001111011000100110001001",
"01010100010000010100011000000000",
"00111110010010000100111001000001",
"10010000100100010000000000100001",
"11110000000000000000000000001101",
"00010000000100010101011000111111",
"11111010101001100011111010001001",
"00001101111110011010101100111110",
"00111111111000000000000000000000",
"11111000010111110011111001010110",
"01000110000000000000010000111101",
"10010001010100110100111101000011",
"00001001100100001001000110010000",
"00000000000000000000110101010101",
"00010001010101100011111111110000",
"11111001100010100011111000010000",
"00001011010100100001000100001111",
"01000010111110010101001000111110",
"00010000000100010000000000011101",
"00111110000100000001000110001001",
"01010001010101101111100000110101",
"01010000000011100001100000001011",
"11110110101100110011111000001100",
"10010001111110100110001100111110",
"11111001011001100011111010010000",
"10010000111111111101100101000000",
"00010001000010101001000100001000",
"10001001000010001000100100010000",
"00000000000001010011110110001001",
"01010011010011110100001101000110",
"11111111101100110011111001001000",
"11110000000000000000000000001101",
"00110010001111100101011000111111",
"00000000000001000011110111111010",
"01010000010110000100010101000110",
"00000000000011010000111000001111",
"00011100011111111111000000000000",
"00100010001010100000111100101100",
"00000000000011000100001000001010",
"00001101000010000001101000001000",
"11111111111000000000000000000000",
"00111101010101100010100001010101",
"00011010000010001001000010010001",
"00100011000000000001010101000110",
"00010111000000111111111101000110",
"10001000000100000010101010010000",
"00001101111101100101010000111110",
"00111111111001100010111001000010",
"11111010001110011110111100001101",
"11110111101111110011111011111110",
"10001001000100010001000000010001",
"11110000000000000000000000001101",
"00111110010101100001110001111111",
"10010000100100011111100111101100",
"11110000000000000000000000001101",
"11010110001111100101011000111111",
"10001001000100000001000111111001",
"10010001111110011101101100111110",
"10001111100011110000100110010000",
"00001111000100000001000101010101",
"00111110000010110101001000010001",
"00100000010000101111100010100011",
"10001001000100000001000100000000",
"10000110001111100001000000010001",
"01010010100100001001000111110111",
"01010001000011100001100000001011",
"00010000001010101001000000001100",
"11110101111111110011111010001000",
"00111110111110011010111100111110",
"11010110010000001111100010110100",
"10010001000010001001000011111111",
"10001001000100000001000100001010",
"00111110100010011000100100001000",
"00000110001111011111100010100100",
"01011000010001010100011000000000",
"00001101001100010100110101010000",
"00111111111100000000000000000000",
"11111000100100100011111001010110",
"00111101111111110101000100111110",
"01001100010001100000000000000011",
"11111111010010000011111001001110",
"00000010011010111011000100001101",
"01010101000101110000110101000000",
"01110001001111101011101110110101",
"00000000000001010011110111111001",
"01010000010011100100110001000110",
"00001111000011110000111100110001",
"11110111001001110011111000001111",
"10010001111101011001101100111110",
"10010000100100010000100110010000",
"00010000000100010101011000001001",
"00001011010100100001000100001111",
"01000010111110000010011000111110",
"00010000000100010000000000100010",
"00111110000100000001000110001001",
"00001011010100101111011100001001",
"00001100010100010000111000011000",
"00111110000110000000111000011010",
"10000010001111101111001000000101",
"11111001001100100011111011110101",
"00110101001111101001000010010001",
"11111111110101000100000011111000",
"00001010100100010000100010010000",
"00001000100010010001000000010001",
"00000100001111011000100110001001",
"01001111010011000100011000000000",
"11111110100000110011111001000111",
"00000000000011011001000010010001",
"01010110001111111111000000000000",
"00111110100010010001000000010001",
"11111010001111101111100100001000",
"00000000000000000000110111111000",
"00111110010101100100000000000000",
"00000100001111011111100011111100",
"01001001010100110100011000000000",
"00111110100100001001000101001110",
"00010000000100011111111110000111",
"11111101111000000011111010001001",
"01000110000000000000010100111101",
"01001000010011100100100101010011",
"11111111000011010000100010010000",
"00011100011111111111111111111111",
"10010000100100011000100000010000",
"00010000000100010101011000001001",
"00000000000000000000000000001101",
"11001001001111100101011001000000",
"00001111000011110000111111111000",
"11110110100001110011111000001111",
"10110010001111100001000000010001",
"01010011000010110101001111111000",
"00000000000000000000110100001011",
"00111110010101100100000000000000",
"10101101001111101111011001110101",
"10011110001111101001000111111000",
"10001000000100000000111111111000",
"00001110000110000000101101010010",
"01110100001111100000110001010001",
"11010000010000100001111111110111",
"10010001000010001001000011111111",
"10001001000100000001000100001010",
"00000111001111011000100100001000"
)
,(
"01001001010100110100011000000000",
"01010011010011110100001101001110",
"00111110111111111000111000111110",
"00000101001111011111100010000000",
"01010001010100110100011000000000",
"11100010001111100101010001010010",
"00001101100100001001000111111101",
"00111111111100000000000000000000",
"00111110000100000001000101010110",
"10010000100100011111100001101000",
"00010001111110000101100000111110",
"00010000000100011000100100010000",
"11110111011000100011111010001001",
"00111101111110000101011100111110",
"01010100010001100000000000000100",
"10010000100100010100111001000001",
"11111000001111110011111000001001",
"11111111000011010000100010010000",
"00011100011111111111111111111111",
"00001111000011111000100000010000",
"10001010000100010010110000100010",
"00111110000100010000101010010001",
"00011010000011111111100000101001",
"00101010000011110011011000100010",
"10001001000100000000101000011100",
"00000000000001010011110100100010",
"01001110010000010101010001000110",
"00000010010001000011111001001000",
"00000001010000100010100100001110",
"11000000000011010010000100000000",
"00000010000001011111111111111111",
"00010000010000100011100000010111",
"00000000001011100100011000000000",
"00000001100001000011111001010101",
"00111110000000010000110100111110",
"00101101010000000000000110111100",
"00011101010000100010100100000000",
"00001000010000001100011000000000",
"01010110001000011000011010001110",
"01000110000010011001000010010001",
"00111110010101100000000000110000",
"10101101100110000000000101100110",
"11110010110000101001111110111000",
"10000101100011111000100111111111",
"00101110010001100101011010001000",
"00111110000110000000111100000000",
"00111110000010000000000101010010",
"01000000010001100000000011011010",
"00011001000011100001111000001000",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"01000110000000000000001000111101",
"11111111100110010011111001111110",
"00111101111011101110011100111110",
"00101110010001100000000000000011",
"00000001110101000011111000101110",
"00111110000000001011010100111110",
"00101110010001100000000011011100",
"00011111001111100101010100000000",
"00000001010110100011111000000001",
"00011110000010000100000001000110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"00000010001111010010001000000100",
"00111110001011100100011000000000",
"10110101001111101111111111010111",
"00000000000001000011110111101110",
"00101110001011100101001101000110",
"00111110000000011010000100111110",
"10101001001111100000000010000010",
"00101010100100000000111000000000",
"00111110010100111000100000010000",
"10010000000010001111000000011011",
"00000000001011100100011000010111",
"00111110000110001000100000010000",
"00011001001111100000000011011110",
"00001000010000000100011000000001",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111101001000100000010000011001",
"01010011010001100000000000000011",
"11111111110010000011111000101110",
"00111101111011100111001100111110",
"01000101010001100000000000000100",
"11000000000011010010111000101110",
"01000110000001011111111111111111",
"00111000001011010000000001000000",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"01000010001010100010110101010011",
"00001010100100010000000000000100",
"00000001000010001000100000010000",
"01000110000000000000001100111101",
"01000000010001100010111001000101",
"10010000000110000000011000001000",
"00001000010000000100011000011000",
"10001000000100000000001100010110",
"00000101000010000100000001000110",
"01010011000000000000110100111101",
"01010000001011010101010001000101",
"01001001010000110100010101010010",
"01001110010011110100100101010011",
"00010000000010000100000011000110",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00001111001000100000010000011001",
"00000100000110010001011000001111",
"00010111000000000011000001000110",
"00010111010101010000111100101100",
"00000100010000100001110000111000",
"11101010010000000001100100000000",
"00001000000001010001000011111111",
"01000000110001100011110110001000",
"00010001000010001001000000001000",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00001111001000100000010000011001",
"00000000001100000100011000000100",
"01010101000011110010110000010111",
"01000010000111000011100000010111",
"00011001100110010000000000100100",
"00001110000110000000111110010000",
"01010110100010000001000000011001",
"01000000000010011001000010010001",
"00010000000011110000000000001001",
"00010000000011110000010000010110",
"10101101100110000000001100010110",
"11110001110000101001111110111000",
"01000000000010011000100111111111",
"00000101000100011111111111001101",
"00111101100010010001000000001000",
"10011110000010000100000011000110",
"11001110100001001001100110001110",
"10011001100110011000111110100000",
"00000100000100011010001010000100",
"00010111000000000010110101000110",
"00010110000100010001011100101100",
"10010000100101101000111110001111",
"10001000000100000001000100001000",
"01000000000010011001000010010001",
"10001110000100000000000000000111",
"10001000000100000000001110000100",
"10011111101110001010110110011000",
"10001001111111111111001111000010",
"10011000100010000000001100010000",
"10000101100110011001100110001111",
"01000101010001100011110110001000",
"11111111001001100011111000000000",
"00000000000001110100001000101001",
"00000000001011010100011000100001",
"01000110000000000000001101000000",
"00010101001111100000000000101011",
"00000000000000010011111011111111",
"11111111111001000000110100111101",
"00111110000000100000010111111111",
"01000010001101011110111100111011",
"11110000001111100000000000000110",
"00000000000000010100000011111111",
"00000000000000010011111000001000",
"00111000001011010100110100111101",
"00000000000001100100001000001010",
"01000000000000000101011101000110",
"00110000010001100000000000000011",
"11100101001111100001011000000000",
"10010001100100000011110111111110",
"00001111111101011111011100111110",
"11111000100101100011111000001111",
"00000000001111100000111100001111",
"00001000100100000000101011111000",
"00010001111101011101110000111110",
"00111110100100010001000110001010",
"10001000000100001111001110100101",
"00111101100010010001000000010001",
"00001000010000000100011001010110",
"01000010001010100000111100000101",
"00101101010001100000000000001001",
"11111110101100100011111000000000",
"00001111111100100000001100111110",
"11110000000000000000000000001101",
"00001000010000100001110001111111",
"00111110000011110000111100000000",
"00000010010000001111101110000010",
"00001101000011100101011000000000",
"00000101111111111111111111100100",
"00010000001010101001000000000010",
"11110001111100110011111010001000",
"01101011001111101001000010010001",
"11110101100111100011111011111011",
"00001010111101111010111000111110",
"00010001000010101001000100010001",
"11111111110000000000110100010000",
"00010111000000100000010111111111",
"00111110111100100010010100111110",
"10001000000100001111010010010000",
"00010001000010101001000100010001",
"11110010000110000011111000010000",
"00101011111111110111111100111110",
"10011001000000000000010001000010",
"00001110000000000000010001000000",
"00010001111111110101111000111110",
"10010000100010100001000110001010",
"00001101001101100000100110010001",
"00000101111111111111111111000000",
"10010001000100010001011000000010",
"10001000000100000001000100001010",
"10010001010101100001100010001001",
"00001111010000000000100110010000",
"00111110100100001001000100000000",
"01001101001111101111010101001100",
"11111111001101010011111011111111",
"10011000100010010001000000010001",
"11000010100111111011100010101101",
"00001001100010011111111111101011",
"10001000000100000000100100001001",
"11111111111111111110010010001101",
"01000000010001101000001000000101",
"00011001000011100001111000001000",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00001111100100011001000000011001",
"00011001000110010000111100001111",
"10000100000101100000100000000101",
"10010111000000000010110111000110",
"00000100000011101001011010101100",
"00101101000000000100000101000110",
"00000110010000100000101000101010",
"00000000001100000100011000000000",
"01000110000000000000001101000000",
"00011010000101110000000000110111",
"00011111001010100001011100010001",
"00011100001101100001000000001110",
"00001000000000000011111101000010",
"01000110000001000000111000011001",
"00101010001011010000000001000001",
"00000000000001100100001000001010",
"01000000000000000011000001000110",
"00110111010001100000000000000011",
"00001110000110000001011100000000",
"01000010001010010001011100010001",
"11010110000010000000000000000101",
"00001010000000000000001001000000",
"00101010001011010100110011010111",
"00000000000001100100001000001010",
"01000000000000000011000001000110",
"00110111010001100000000000000011",
"00000011000011110001011000000000",
"01000000100110011000100000010000",
"00001010100010011111111110111010",
"01000110000000000000100001000010",
"00111110010101100000000000110001",
"00111101000110001111111000100010",
"01000110000010000100000001000110",
"01000110000101100000000100000000",
"00111101000000010101101010001100",
"00000010010110101000110001000110",
"10001100010001100000111000011001",
"00111101000000110000000101011010",
"00100011001111000000000000000010",
"00000000000001100100001000101010",
"00111110000000000010110101000110",
"00000100001111011111111111100110",
"01001100010011110100100000000000",
"11111111111001000000110101000100",
"00111110000000100000010111111111",
"00001000100100001110110011000111",
"00010000000100010000101010010001",
"00101010001011010100110010001001",
"00001000000000000000011101000010",
"01000000000000000011000001000110",
"01000110000101110000000000000100",
"00111110000101100000000001000001",
"00000100001111011111111110111010",
"01000111010010010101001100000000",
"11111111110100010011111001001110",
"00101100001000100000111100001111",
"00111101111111111111011001000010",
"00001001001000110000000000000001",
"00000010010110101000110001000110",
"01000110000010000100000001000110",
"00001111000101100000000100000000",
"00000000000000100011110100010111",
"10010001100100000101001100100011",
"11111111100000000011111000001001",
"00010001111111111101011000111110",
"00111110111111111001010100111110",
"00010000000010101111111111011101",
"01010110001000010001011110001001",
"01000000000010011001000010010001",
"00100000010001100000000000000111",
"11111111011100000011111000000000",
"10011111101110001010110110011000",
"10001001111111111111001111000010",
"00100011000000000000001000111101",
"00001001100100011001000000111110",
"10001001000100010001000001010110",
"00111101000000000111111000111110",
"00111110111111111111001000111110",
"00000100001111011110101100011000",
"00101110001011100101010100000000",
"11101111001111100101011001010010",
"00000000000000110011110111111111",
"10010000010100100010111001010101",
"00010111000011100000100010010001",
"00000001010000100010100100010000",
"00010000000100010010000100000000",
"11111111100111100011111010001001",
"10000110001111100000111001010110",
"00000000000000100011110111111111",
"11100010001111100010111001010101",
"11101010111001100011111011111111",
"00101110000000000000001100111101",
"00111110010101100101001000101110",
"00000010001111011111111111110000",
"01010110010100100010111000000000",
"00111101000000000010010100111110",
"10010000001011100000000000000001",
"00101010000011111001000100001000",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00111110100010010001000000010001",
"00001110010101101111111101100000",
"00111101111111110100100000111110",
"00101110010001000000000000000010",
"00111110111111111101110000111110",
"00000100001111011110101010101000",
"00101110001011100100010000000000",
"01000101001111100101011001010010",
"00111110000011100101011011111111",
"00000011001111011111111100101101",
"01010010001011100100010000000000",
"11101001110010010011111001000011",
"11011000010001100000111001000100",
"00000101001111010000000111111111",
"00101110010001000101010100000000",
"01000110010000110101001000101110",
"01000110000000101111111111101100",
"01000110000111000000000000010010",
"00101100000101110000000000010010",
"01000110000000011011111101000010",
"00001110000000101111111111100000",
"00010111000000010000000001000110",
"11000110000110000000111000101010",
"00000010000100000000101001010100",
"00000001100010000001000000010110",
"00000100000010100100110001000110",
"01000110010101100001110000101100",
"01000010000000110000101001001100",
"11000110000011100000000101010111",
"01000110000000000000000100000000",
"00101100001011010000000011111111",
"00000000000011000100001000001010",
"11011000010001100000111000001000",
"10101011001111100000000111111111",
"00000001001111000100000011011010",
"00000000111111100100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000010010100101000000",
"00101101000000001111110101000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000100010110",
"00101100001011010000000011111100",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"00000011010000000001000000000001",
"11111011010001100000000000000001",
"00001010001011000010110100000000",
"00001000000000000000111101000010",
"11111111110110000100011000001110",
"00001110010001100000110100000001",
"01000000101111010000010000000000",
"01000110000000000000000011101010",
"00101100001011010000000011111010",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"11010111010000000001000000000001",
"11111001010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000000110001000100000000010000",
"00000000111110000100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000001011000101000000",
"00101101000000001111011101000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000010011110",
"00101100001011010000000011110110",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"10001011010000000001000000000001",
"11110101010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000000011110000100000000010000",
"00000000111101000100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000000110010101000000",
"00101101000000001111001101000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000001010010",
"00101100001011010000000000011011",
"00000000000010010100001000001010",
"00001010010011000100011000001000",
"00111111010000000001000000000011",
"00011010010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000111001000010",
"00000011000010100100110101000110",
"00001010010011100100011001010110",
"00100111010000000001000000000011",
"00011001010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000111001000010",
"00000011000010100100110101000110",
"00001010010011100100011001010110",
"00001111010000000001000000000011",
"01000110000011100000100000000000",
"00101010000101110000000000010000",
"01000110000000000000010101000010",
"00010000000000110000101001001110",
"00000000010001100000111010001000",
"01000010001010100001011100000001",
"01001110010001100000000000111000",
"00011010000110100000010000001010",
"01000000010001100001101000011010",
"00011101100100000001011000001001",
"10011101100111011000111000000010",
"00000010000100001001110110001110",
"00011010010000100101110000101101",
"00010000000110000000111000000000",
"00000010000100000000000110001000",
"00011111010111000010110100010110",
"00010111000000000000001101000010",
"00010001000010100000111000100001",
"10001110000000110001011000000010",
"10001001000011100000111000001110",
"01000000000010000000100110001000",
"01000110000011101111111000110001",
"01000100000000011111111111011000",
"11111111110101001100011000111101",
"11111111111011000100011010000010",
"00101100000111000101000100000010",
"10010000111111111111011001000010",
"10010111110011100000100110010001",
"00000000000100001100011010101100",
"01010100000000001101011010011100",
"01000010000010100010110000101101",
"10011110000010000000000000000101",
"00000000000000000000111001000000",
"00001010001011000010110101010101",
"00001000000000000000010101000010",
"00000000000000010100000010011000",
"00000000110100101010001000001000",
"00001010001011000010110101010010",
"00001000000000000000011001000010",
"00001110010000001001011110001110",
"00101101010100110000000000000000",
"00000101010000100000101000101100",
"01000000100110100000100000000000",
"10100010000010000000000000000001",
"10000001111111111110010011000110",
"00010110000100000000001001011010",
"00111110000110101000100000010000",
"11101000010001101110101001000010",
"11010100110001100000000111111111",
"11000110001111011000000111111111",
"00010000100000101111111111100100",
"01010110000000000001110001001010",
"01000010000010100010110000101101",
"01010010000010000000000000000101",
"00000000000000000000111101000000",
"00001010001011000010110101001110",
"00001000000000000000010101000010",
"00000000000000100100000001010011",
"01010011000100000101010000001000",
"00101101010101000000000000011100",
"00000101010000100000101000101100",
"01000000010101000000100000000000",
"01010101000000000000000000001111",
"01000010000010100010110000101101",
"01010101000010000000000000000101",
"00001000000000000000001001000000",
"00010000110001100100111101010110",
"00000001110000101001110000000000",
"00000010010110100001100000000000",
"10000010111111111110100011000110",
"10001000000100000001011000010000",
"11101001111000000011111000011010",
"01010011000000000000011000111101",
"01001001010100110101010001000101",
"10100100001111100100111101001111",
"00000100100100000000100100001000",
"10011000000001000001000010011000",
"00010000100110000000010000010000",
"00000100000100001001100000000100",
"10011000001000100010000001001110",
"00010000010001100000010000010000",
"10011000001000100010000000000000"
)
,(
"01000110000001001000100000010000",
"00100010001000000000000000011000",
"00111101111111110000101000111110",
"01000101010001110000000000000110",
"01001111010010010101001101010100",
"00111110000000000001000001000110",
"01011010010101011110011100111010",
"00001001010011000100011000000001",
"00000100000000000100011000000010",
"00111110000011100001011100001111",
"01011010010101001110011101100110",
"00111110001000110100111000000001",
"01011010010100101110011101011110",
"01010111001111100101011000000001",
"00000001010110100100111011100111",
"00111110000000000001101001000110",
"00010000010001101110011100010010",
"00111101000000010101101000000000",
"00000010000010010100110001000110",
"00000000001100000100001000101100",
"00111110000000000001000001000110",
"00000000010001101110011011111110",
"00110011001111100000111000000100",
"00111110001000110100111011100111",
"00111110010101111110011100101110",
"00011010010001101110011100101010",
"11100110111010000011111000000000",
"00000010111111111101010001000110",
"11111111110101000100011001010101",
"00001001010011000100011000000001",
"11111111111110010100001000000010",
"00000001111111111101010001000110",
"00000010111111111101010001000110",
"00000010000010010100000001000110",
"00000010000010010100100001000110",
"01001100010001100000010000010110",
"00010111010101010000001000001001",
"01001100010001100010010101010110",
"01001000010001100000000100001001",
"01000110000110000000001000001001",
"01000110000111000000001111111111",
"10010001000000010000100101001000",
"01000110100010000001000000001010",
"00111101000000011111111111010100",
"01000101010010110000000000000100",
"00101101000011100011111101011001",
"00000000000001110100001000101100",
"11111111100010000011111000001000",
"10001101111111111111010001000000",
"00000101111111111111111111111100",
"11011010100101101101001110000010",
"00101101100111101000111010011100",
"00000000000010010100001000110110",
"00111110100110000000001100010000",
"11110010010000001111111101101110",
"10010111100011110000100111111111",
"10000101100011111001100110011001",
"00000011001111011000100000010000",
"01011001010001010100101100000000",
"00011110111111111100011100111110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"00000100001111010010001000000100",
"01010010010011110101011100000000",
"11010100110001100000100001000100",
"01001000010001101000001011111111",
"01001100010001100000000100001001",
"11010100110001100000000100001001",
"00000101001111011000000111111111",
"01010010010000010101000000000000",
"11010100110001100100010101010011",
"01001100010001101000001011111111",
"01001000010001100000001000001001",
"11000110010101010000001000001001",
"00111101100000011111111111010100",
"01000101010100100000000000001101",
"01010010010011110101010001010011",
"01001110010010010010110101000101",
"01010110010101000101010101010000",
"00111110000110000000111000001110",
"00001010001111011111111110111111",
"01010110010000010101001100000000",
"01001110010010010010110101000101",
"00111110010101000101010101010000",
"10111111001111101111111111101001",
"00000000000001010011110111111110",
"01010010010001010101010101010001",
"11010110000010001001000001011001",
"00001110111111101110010100111110",
"11100110011001000011111010010000",
"11001100000110000000001100001111",
"00000101110000101010110010010111",
"01000000100011101000101000000000",
"10101101100110000000000000000001",
"11100011110000101001111110111000",
"10001001000100010000100011111111",
"01010010000000000000011000111101",
"01001100010010010100011001000101",
"11111111110100010011111001001100",
"11111111111111111111000000001101",
"00000110001111010000000100000101",
"01000011010000110100000100000000",
"10010000010101000101000001000101",
"00000010000011101001000000001000",
"00000010000011100001110100010110",
"00111000001011010001110100010110",
"10010000000000000100001101000010",
"00011000000011100000001010011101",
"00010001000000000000111001000010",
"00011101000100000001000100010110",
"00111110000000101000100000010000",
"00101010010000000000000000111011",
"00111110000100000000100000000000",
"10001110100111101110001101001011",
"10100000110011101000010010011001",
"10000100100110011001100110001111",
"10010110110100111001011010100010",
"00001001010000101001110011011010",
"00010000000100010000111000000000",
"00111110100100010001000110001000",
"00010000000010000000000001001100",
"00011000000000101000100000010000",
"01000000000101100001101000011010",
"10001001000010011111111110111000",
"01000101000000000000011000111101",
"01000011010001010101000001011000",
"10010000100100010101011001010100",
"00000000001001000100000000001001",
"10010001000000101001110110010000",
"00000011100100001001000100010110",
"10011000001000110100111000010001",
"01000110000100010000001100010000",
"10011000001000110000000000010000",
"01000110000100010000001100010000",
"10011000001000110000000000011000",
"10001001000100010000001100010000",
"10011000100010010001000100010000",
"11000010100111111011100010101101",
"00001010100010011111111111010110",
"00001000100100000011110100001010",
"10011001000100001000001010010000",
"00011101000000001001101001000010",
"00011000000011100000001000001110",
"11111111000011010000111100110110",
"00011100011111111111111111111111",
"00011111001010100001011100010001",
"00000000100000010100001000011100",
"00010110000011110000101010010001",
"00100011010101010001101010010000",
"11000110100001001001000000011001",
"00010001100111000000000010000000",
"10101010000010001001000010001010",
"01001001000000000011000011000010",
"00000010000111010000101101010011",
"00011100000000001111111101000110",
"00101100001011010101001100000000",
"00000000000010000100001000001010",
"00111111010001100000100000001000",
"00000000000011110100000000000000",
"00101100001011010101001000000000",
"00000000000001010100001000001010",
"00000010010000001001111000001000",
"00010000100110000000100000000000",
"00011100000000001000000001000110",
"00011000000000110000111100100010",
"00011101000111010000101101010100",
"00000001010000100100001110011011",
"10010001100100000000001000000000",
"00000011000100000001000100001001",
"10011000001000110100111000010001",
"01000110000100010000001100010000",
"10011000001000110000000000010000",
"01000110000100010000001100010000",
"10011000001000110000000000011000",
"00010001100010100000001100010000",
"00000101010000100001110001010101",
"00010000000110100001000100000000",
"01010111100010010000001100011000",
"10001000000100000000000100010000",
"01100001010000000000100000001110",
"10001001000010010000100011111111",
"01010110000000100000111000111101",
"01000000000010011001000010010001",
"10010000000111010000000000011010",
"11111111000011010001100000000010",
"00011100011111111111111111111111",
"00001010000111110011100000101101",
"00000000000001000100001000001110",
"00111101100010011000100000001010",
"10011000100010000001000000001000",
"11000010100111111011100010101101",
"00001001100010011111111111100000",
"10010000100100010011110101010110",
"00000010000011101001000000001001",
"00000010000011100001110100010110",
"00111000001011010001110100010110",
"10010000000000001000001001000010",
"10101100100101111101011110000010",
"00000000011100001100001000011101",
"00011001000011100001111000001110",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"01011010000101100101001100010110",
"00010001100010000001000000011100",
"00111110000011110000101010010001",
"01010010010000101111111110011111",
"00001110000111100000111100000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11100100011101100011111000100010",
"00000000001010111001101000001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110111001000110001100111110",
"00101010000100011110010010110101",
"01000111000000000010001101000010",
"01000110111000111110110100111110",
"00100011001111100000000000011000",
"10111011001111100001000011100100",
"10010111100100011001000000000101",
"00011000000000100000111100001111",
"10001000000100000001101000011010",
"11100100001001100011111000010110",
"00111110000000000001101001000110",
"10001000000100001110001111001110",
"00001010000010001001000010011000",
"00011010000110000000001000001110",
"01111001010000000001011000011010",
"00010000100010000000100111111111",
"00000000000010100011110110001001",
"01100100011011100111010100100000",
"01101110011010010110011001100101",
"10111101010001010110010001100101",
"11111111111111111100110000001101",
"01000110000011100000001000000101",
"00011001000000100000101001110100",
"00010000000010101001000100010110",
"00000010000011100000111010001000",
"10010000000111010001011000011101",
"00010000000011110000111100001000",
"11010010001111100001011100001111",
"00010111000011110001000011111101",
"11111111001100100011111001010110",
"00000000010100000100001000101011",
"00111110100010000001000000001000",
"00101100000001111111111111001100",
"00001101000000000010011001000010",
"00000101111111111111111111001100",
"01110100010001100000111000000010",
"00010110000110010000001000001010",
"10001000000100000000101010010001",
"00011010010101010000111100001111",
"11111101101000110011111000011010",
"01000110000110100001101001010101",
"00111110000000100000101001111000",
"00011100010000001111111100000000",
"11100100000010110011111000000000",
"00000000001011000010011000001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110111000111010001100111110",
"00100101001111101110001111110101",
"00000000000000010100000011100010",
"00000000010011110011110110001000",
"00101010001010100010101000101010",
"00101010001010100010101000101010",
"01110100011000010110010000100000",
"01110100011100110010000001100001",
"00100000011010110110001101100001",
"01110010011100100110111101100011",
"01100101011101000111000001110101",
"01101000011101000010000001100100",
"01100111011101010110111101110010",
"01101110011010010010000001101000",
"01100001011010010111010001101001",
"01101111011000110010000001101100",
"00100000001011000110010101100100",
"01100011011100100110111101100110",
"01100001001000000111001101100101",
"01110011011001010111001000100000",
"01110100011100100110000101110100",
"00101010001000000010000100100000",
"00101010001010100010101000101010",
"00001101001010100010101000101010",
"00000101111111111111111111001100",
"00001010011111000100011000000010",
"01111000010001100010110000000010",
"00100010001011000000001000001010",
"00001101000000000000111101000010",
"00000101111111111111111111111100",
"00001010011011000100011000000010",
"01111100010001100000111000000001",
"01000110010101100000000100001010",
"01010111000000010000101001010100",
"00000011000010100100111101000110",
"00000000111100000100011001010111",
"01000110000000111010000100111110",
"00100010000000100000101001010100",
"00001010011101000100011000001111",
"01110000010001100000111000000001",
"00101100000010100000000100001010",
"00001101000000000100101101000010",
"00000101111111111111111111001100",
"00010000010100011001000000000010",
"11011111011100000011111000011101",
"00111000111111101101100100111110",
"01000110000100010001111110010000",
"00011001000000100000101001110100",
"01000010000111000000010000010110",
"00001110000100010000000000001111",
"00011101000101100000001010001001",
"11111111111111111100110000001101",
"00011101010000000000000100000101",
"00001010011100001100011000000000",
"00001010011011000100011010000001",
"11111111111111000000110100000010",
"10001000000000010000010111111111",
"00001010011111000100011001010110",
"00111110000111010000001000001110",
"01011111001111101110000000001011",
"00111110010001110000000111100000",
"00010100010001101110001001000110",
"11100010011111000011111000000000",
"00000010000010100101010001000110",
"01000110000001000001000100111110",
"00110110000000100000101001110000",
"00010110000000000001101001000110",
"01010110111000100010110100111110",
"00000011000010100100111101000110",
"01011000001111100101011100111101",
"01000010001011001001000000000011",
"00010110100100010000000001100001",
"00111000001011011000100000010000",
"10010000000000000101100001000010",
"00011110000011100001110110000010",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"01010011000101100010001000000100",
"00001111000111000101101000010110",
"01000010110111111011101000111110",
"00010001100100010000000000001011",
"00111110010100101000100100010000",
"00101000010000001111110011001100",
"10011000100010000000100000000000",
"00011001000011100001111000001111",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00001101111000100100011100111110",
"00000100000000000010110111010010",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"10000110001111101110001000110100",
"00000010000011100000101011100010",
"00010110000110100001101000011000",
"00001001111111111010001101000000",
"00001010011111000100011001010110",
"00000000000100111100001010110101",
"00000010000010100110110001000110",
"11111111111111111111110000001101",
"00000010000011100000000100000101",
"11011111011000010011111000011101",
"00000001110111111011010100111110",
"11100001100111000011111001000111",
"00111110000000000001010001000110",
"10001000000100001110000111010010",
"00000011011010000011111000001110",
"00000000000110100100011000110110",
"11010100010001100101010100010110",
"10000011001111100000000111111111",
"00000000000010110011110111100001",
"01110010011011100111010100100000",
"01101100011011110111001101100101",
"01001110011001000110010101110110",
"00111101001000100101010100111101",
"01001001010001000000000000000011",
"00000011001111010101001001010010",
"01001110010010010100001000000000",
"00000000000000110011110101010100",
"01010000010011110010111101010111",
"01010010000000000000001100111101",
"11010100010001100100111100101111",
"00001110010101100000001011111111",
"00000011000010100100110101000110",
"00000001000010100101010001000110",
"00000001111111111101010001000110",
"00000100000010100100110101000110",
"11111111111110000100001000110110",
"00000010111111111101010001000110",
"00000100000010100100110101000110",
"00010111000000000001101001000110",
"00001010010101000100011000100001",
"00001110010101100001011000000010",
"00000011000010100100110101000110",
"00000001000010100101010001000110",
"11111111110101000100011000001111",
"00000011001111010000101000000001",
"01010111001011110101001000000000",
"10010000100100010101010101001000",
"00001010010100000100011000001001",
"00100000000100000101010100000010",
"00101100000111000000111100001111",
"00100010000000000000100001000010",
"00000001000010100101000001000110",
"00001001001111011000100100010000",
"10011111101110001010110110011000",
"10001001111111111110001011000010",
"11010100110001100011110101010111",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01000111111000001110000100111110",
"10010000111000010001100100111110",
"01000110111000010001010100111110",
"11010011001111100000000000011010",
"11111111011110100011111011100000",
"00000000000100110100001000101011",
"10011011100110111001101110011011",
"00011111001000000001000001010101",
"01010000110001100010001001010101",
"00011100000000100001000000001010",
"10001000100010000000000100010000",
"10000001111111111101010011000110",
"11111111110101001100011000111101",
"11010100010001100101010110000010",
"00001000100100000000000111111111",
"00011010111111111001000100111110",
"00100010000110100001101000011010",
"00011101010000100001111100101001",
"00111110010001111001000000000000",
"00111110000100011110000010010110",
"11001011001111101110000011001110",
"11100000110111100011111011100000",
"00111110000000000001101001000110",
"10001001000100001110000010000110",
"01000000111111110010101100111110",
"00001010100010000000000000000100",
"11010100110001100000111000001010",
"00001010001111011000000111111111",
"01001111010011000100001100000000",
"01000110001011010100010101010011",
"00111110010001010100110001001001",
"01010101001000101111111011111011",
"00111101111111111010111000111110",
"11111111101010010011111001010110",
"01000011000000000000101100111101",
"01010100010000010100010101010010",
"01001001010001100010110101000101",
"11010100110001100100010101001100",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01001000111000000100000100111110",
"00111110111000000111100100111110",
"00011010010001101110000010001100",
"11100000001101000011111000000000",
"11000110111111101101101100111110",
"00111101100000011111111111010100",
"01010000010011110000000000001001",
"01000110001011010100111001000101",
"11000110010001010100110001001001",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11100000000101000011111001000111",
"11100000010011000011111001010000",
"01000110111000000100100100111110",
"00000111001111100000000000011010",
"11111111111111000000110111100000",
"01010011000000100000010111111111",
"01001110000111000101101000010110",
"00111110000000001111000001000110",
"00111110000010000000000010111110",
"00001000100100001111111010011100",
"11111111111111111111110000001101",
"00010110010100110000001000000101",
"00011101100100000001110001011010",
"00000010100010000001000000000010",
"11010100110001101000100000010000",
"00001011001111011000000111111111",
"01001100010001010100010000000000",
"00101101010001010101010001000101",
"01000101010011000100100101000110",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"10111111001111100100011100000001",
"11110111001111100100111011011111",
"11011111111101000011111011011111",
"00111110000000000001101001000110",
"11111100000011011101111110110010",
"00000010000001011111111111111111",
"00011100010110100001011001010011",
"00000000111100000100011001001110",
"00001000000000000110100100111110",
"10010000111111100100011100111110",
"11111111111111000000110100001000",
"01010011000000100000010111111111",
"10010000000111000101101000010110",
"10001000000100000000001000011101",
"11000110100010000001000000000010",
"00111101100000011111111111010100",
"01001001010001100000000000001101",
"01010000001011010100010101001100",
"01010100010010010101001101001111",
"00001000010011100100111101001001",
"01000110000000000000100100111101",
"00101101010001010100110001001001",
"01000101010110100100100101010011",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"01011011001111100100011100000001",
"10010011001111100100110011011111",
"11011111101001100011111011011111"
)
,(
"00111110000000000001101001000110",
"11110101001111101101111101001110",
"11111111110101001100011011111101",
"00000000000011000011110110000001",
"01001100010000110100111001001001",
"00101101010001010100010001010101",
"01000101010011000100100101000110",
"11110000010001101001000010010001",
"01000000010001100001110000000000",
"00011101100100000001011000001001",
"10011101000000010001000000000001",
"00001111000100000101011010011101",
"00000001000000010001000010011101",
"00111101100010011000100000010000",
"01001110010010010000000000001000",
"01000100010101010100110001000011",
"00011100010001110100010001000101",
"01000000010001100001101000011010",
"00111101000000100001011000001001",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"00111110100100001001000100000001",
"00001000100100001111111111000010",
"11011110111101000011111001000111",
"11011111001011000011111001010100",
"00100111001111101000101000010001",
"00111110100010100001000111011111",
"00011010010001100000000010111110",
"11011110111000000011111000000000",
"10010000111111011000011100111110",
"00010000000000100001000100001000",
"11111111110101001100011010001001",
"00000000000001010011110110000001",
"01000011010011110100110001000010",
"11111111110101001100011001001011",
"00001101000010001001000010000010",
"00000101111111111111111111111100",
"01011010000101100101001100000010",
"11110000010001100001000000011100",
"11111111011111000011111000000000",
"00111110010001110000100010010000",
"00010110010001101101111010101110",
"11011110111001000011111000000000",
"00111110000000001111000001000110",
"10001010000100011101111011011110",
"01010101000000000111010100111110",
"00000001111111111101010001000110",
"00111110000000000001101001000110",
"00111001001111101101111010010010",
"00001101000010001001000011111101",
"00000101111111111111111111111100",
"01011010000101100101001100000010",
"00010000000000100001000100011100",
"11111111110101001100011010001001",
"00000000000010010011110110000001",
"01000100010000010100010101010010",
"01001100010010010100011000101101",
"11111111110101001100011001000101",
"11010100010001100101010110000010",
"10010000100100010000000111111111",
"00011100000000001111000001000110",
"00010110000010010100000001000110",
"00010000000000010001110110010000",
"01010110100111011001110100000001",
"00010000100111010000111100010000",
"10001000000100000000000100000001",
"11011110010010000011111001000111",
"11011110100000000011111001010011",
"11011110011111000011111000010000",
"00000000000101000011111000010001",
"00111110000000000001101001000110",
"00111110100010011101111000110110",
"00001000100100001111110011011100",
"11000110100010000001000000000010",
"00111101100000011111111111010100",
"11011110011000000011111000001110",
"00111110000011100010001101001110",
"00100011010011101101111001011010",
"11011110010101000011111000001110",
"01001111001111100010001101001110",
"00000000000010010011110111011110",
"01000100010000010100010101010010",
"01001110010010010100110000101101",
"11111111110111000011111001000101",
"00111101111111111101100100111110",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"11110011001111100100011100000001",
"00101011001111100100111111011101",
"11011110001010000011111011011110",
"01000110111111111110001000111110",
"11100011001111100000000000011010",
"11111100100010100011111011011101",
"10000001111111111101010011000110",
"11111111110101001100011000111101",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010011011101110111001110",
"00000011001111101101111000000110",
"11111111101111010011111011011110",
"00111110000000000001101001000110",
"01100101001111101101110110111110",
"11111111110101001100011011111100",
"00000000000011110011110110000001",
"01001111010100000100010101010010",
"01001001010101000100100101010011",
"01000110001011010100111001001111",
"11000110010001010100110001001001",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011101100110000011111001000111",
"00111110000000000001001001000110",
"11100001001111101101110111001110",
"11111111100001010011111011011101",
"00111110000000000001101001000110",
"00101101001111101101110110000110",
"11111111110101001100011011111100",
"00000000000010110011110110000001",
"01001001010100110100010101010010",
"01000110001011010100010101011010",
"11000110010001010100110001001001",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"00011011000110110001101100011011",
"00111110110111010110000100111110",
"00011010010001101101110110110000",
"11011101010110000011111000000000",
"10000001111111111101010011000110",
"00000000000011000011110101010110",
"00101101010101000100010101010011",
"01000101010011000100100101000110",
"01000101010101000100000101000100",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"00011011000110110001101100000001",
"11011101001101000011111000011011",
"01001001110111011000001100111110",
"01001100110111010110100100111110",
"01000110110111010110010100111110",
"00100011001111100000000000011010",
"11111111110101001100011011011101",
"00001010001111010101011010000001",
"01001001010100100101011100000000",
"01000110001011010100010101010100",
"11000110010001010100110001001001",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011101000001000011111001000111",
"11011101001111000011111001001010",
"01000110110111010100111100111110",
"11110111001111100000000000011010",
"11111111111111000000110111011100",
"01010011000000100000010111111111",
"01010010000111000101101000010110",
"00111110000000001111000001000110",
"00111110000010001111110110101110",
"00001000100100001111101110001100",
"11111111111111111111110000001101",
"00010110010100110000001000000101",
"00010000000000100001110001011010",
"11111111110101001100011010001000",
"00000000000010100011110110000001",
"01010100010010010101001001010111",
"01001001010011000010110101000101",
"11010100110001100100010101001110",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01000110110111001011010100111110",
"11101011001111100000000000010011",
"11011100111111100011111011011100",
"00111110000000000001101001000110",
"11111100000011011101110010100110",
"00000010000001011111111111111111",
"00011100010110100001011001010011",
"00000000111100000100011001001110",
"00001000111111010101110100111110",
"10010000111110110011101100111110",
"11111111111111001000110100001000",
"11010011100000100000010111111111",
"00010000100111001101101010010110",
"00000010000100000000001000011101",
"11010100110001101000100100010001",
"00001011001111011000000111111111",
"01001100010010010100011000000000",
"01010100010100110010110101000101",
"01010011010101010101010001000001",
"00001100001111010101011000001000",
"01010100010001010100011100000000",
"01001100010010010100011000101101",
"01010100010000010100010001000101",
"11111111110101001100011001000101",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010010011101110001001110",
"10010000100100011101110010000110",
"01111111001111100000111000001001",
"00100011010011100000111011011100",
"00111110110111000111100100111110",
"00010000000100011101110010001100",
"01101111001111100000111010001001",
"00100011010011100000111011011100",
"00111110110111000110100100111110",
"00011010010001101101110001111100",
"11011100001001000011111000000000",
"11000110111110101100101100111110",
"00111101100000011111111111010100",
"01001100010001100000000000001010",
"00101101010010000101001101010101",
"01000101010011000100100101000110",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"00000011001111100100011100000001",
"11011100001111000011111011011100",
"11011100001110000011111000001110",
"00111110001000110100111000001110",
"01000101001111101101110000110010",
"11110000010001101001000111011100",
"11111100101101000011111000000000",
"00011010010001100000100010010000",
"11011011111001000011111000000000",
"00010001111110101000101100111110",
"00010001000010101001000110001010",
"11000110100010010001000000000010",
"00111101100000011111111111010100",
"01000101010100100000000000001011",
"01000101010011010100000101001110",
"01001100010010010100011000101101",
"00000000000100000100011001000101",
"00111101111111111011000100111110",
"00111110000000000001000101000110",
"00001101001111011111111110101010",
"01010011010000100100000100000000",
"01010100010101010100110001001111",
"01001001010001100010110101000101",
"11010100110001100100010101001100",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01010010110110111001110100111110",
"00001101110110111101010100111110",
"00000110000000000000000000000000",
"11111111111111111101100000001101",
"10010000100100010000001000000101",
"00000000001001010100000000001001",
"00011110000011100000001000010000",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"00001010000111100010001000000100",
"00010000110110111100011100111110",
"00111110010100100000111000011101",
"01010010000111011101101111000000",
"01010011110110111011101100111110",
"00001000100100000001101000011010",
"10011111101110001010110110010110",
"10001001111111111101010111000010",
"00111110000000000001101001000110",
"11010100110001101101101101010110",
"00001100001111011000000111111111",
"01010100010011100100010100000000",
"01010011010001010100100101010010",
"01001100010010010100011000101101",
"11111111110101001100011001000101",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010010111101101100110110",
"00011010010001101101101101101110",
"11011011001011000011111000000000",
"10000001111111111101010011000110",
"01010010000000000000111000111101",
"01000100010001000100000101000101",
"01001001010101000100001101001001",
"01010010010000010100111001001111",
"11111111110101001100011001011001",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010100011101101100001010",
"00111111001111101101101101000010",
"11011011001111000011111011011011",
"00111110000000000001101001000110",
"11010100110001101101101011111010",
"00000100001111011000000111111111",
"01000111010000010101000000000000",
"11111111110101001100011001000101",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00010111010001101101101011100010",
"11011011000110000011111000000000",
"01000110110110110001010100111110",
"11010011001111100000000000011010",
"11111111110101001100011011011010",
"00000000000001010011110110000001",
"01011000001011010101010001000001",
"11110111001111100000111101011001",
"00000000001001000100001000001000",
"00001100010000100011010100001111",
"01000110000000100001110100000000",
"00000010000101100000000000010000",
"11010111111100000011111000001111",
"00000000000011000100001000110110",
"00000010000111010000100010010000",
"00010000000000100001011001010110",
"11111111111000000100000010001000",
"00000000000000100100000000001000",
"00001101001111010101011000001001",
"01000001010010000100001100000000",
"01000011010001010100011101001110",
"01010011010100100100000101001000",
"00111110000011110101010001000101",
"00100000010000100000100010111010",
"00110101000011100000111100000000",
"00001000000000000000011001000010",
"00000000001001000011111000001111",
"00000000000011000100001000101011",
"00000010000111010000100110010001",
"00010000000000100001011001001110",
"11111111111001010100000010001000",
"00000010010000000000101000001010",
"00111101010101100000100100000000",
"01001110010010010000000000001010",
"01001110010000010101010001010011",
"01000110010011110100010101000011",
"10001000001111100000111100001111",
"00100101010000100010101111111111",
"00110101000011110000100000000000",
"00011101000000000000110001000010",
"00000000000100000100011000000010",
"00111110000011110000001000010110",
"01000010001101101101011101111010",
"00001000100100000000000000001100",
"00010110010100100000001000011101",
"01000000100010000001000000000010",
"01000000000010001111111111100000",
"00001010000010100000000000000010",
"01000011000000000000011000111101",
"01010100010101000101001101000001",
"10010000000010001001000001001111",
"00000000000101010100001000110101",
"00010000000011110000001010011101",
"00011100000100010010010000000010",
"00011100001101100000111100110110",
"00011001000000000000011001000010",
"11101101010000001001110110011101",
"01000010000011100000101011111111",
"00010000000010000000000000000100",
"00111101100010010000001000011101",
"10001000000100000000111010010001",
"11111111110100010011111001011010",
"00000000000000110100001000110101",
"00001000101111010000101000001010",
"00000000001101011101110100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110110110100011101100111110",
"11010001000011011110111101011000",
"00011110000001000000000000110101",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"00100101001111100010001000000100",
"01000110000000100001110111011010",
"00000010000101100000000000010000",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"11000101000011011101101000010000",
"00011110000001000000000000110101",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"11111101001111100010001000000100",
"11011000100000100011111011011001",
"00100000000000000000101000111101",
"00100000011101000110111101101110",
"01101110011101010110111101100110",
"00100000000000000000101001100100",
"01100011001000000110011001101111",
"01110011011100110110000101101100",
"01100011000000000000110000100000",
"01110100011100110110111001101111",
"01110100011000110111010101110010",
"10010000001000000111001001101111",
"10001010000100011001000100001000",
"10010000000000000001110101000010",
"10001111001111100000111000001000",
"00001111001101010001110000000111",
"00010110010100100000001000011101",
"00110110000011110000111100000010",
"00000000000001010100001000011100",
"11101101010000000000101000001010",
"10001000000100000000100111111111",
"00000111011101000011111000001111",
"00000000010110010100001000011111",
"00000000001101110011101100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110110110011001001100111110",
"00011001000011011110111010110000",
"00011110000001000000000000110111",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"01111101001111100010001000000100",
"10011001001111100001000011011001",
"00110101110100010000110111101110",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11011001011001100011111000100010",
"01000110000000100001110100010000",
"00000010000101100000000000010000",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"11010101001111101101100101010000",
"00010011001111100000111111010111",
"00000000001100010100001000000111",
"01000010001101011101101000001111",
"00001111000011110000000000011110",
"00010110010010100000001000011101",
"10110000001111100001000000000010",
"00000101010000100011010111111110",
"00001010000010101000100100000000",
"00011101000010001011110100001010",
"00000010000101100101011000000010",
"11111111110111100100000010011011",
"00011101000010001001000000001000",
"00000010000101100100111000000010",
"11001000010000001000100100010000",
"00110111001110110000110111111111",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11011001000000100011111000100010",
"00001101111011100001111100111110",
"00000100000000000011010111010001",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"00011101000100001101100011101100",
"00000000000100000100011000000010",
"00001110000111100000001000010110",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11011000110101100011111000100010",
"00000000001101110000010000001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00010000110110001100001100111110",
"11101101110111100011111010001000",
"00111101110101110100001100111110",
"01101110001000000000000000010011",
"01100110001000000111010001101111",
"01100100011011100111010101101111",
"01100001011010000010000000101100",
"01100101011011000110010001101110",
"00100000000000000010000000100000",
"01110101001000000110011001101111",
"01100110011001010110010001101110",
"01100100011001010110111001101001",
"01101010011000100110111100100000",
"00100000011101000110001101100101",
"01100001001000000111010001100001",
"01100101011100100110010001100100",
"00000111001000000111001101110011",
"01110100011001010110110100000000",
"00100000011001000110111101101000",
"01011000010001010000000000001011",
"01010100010101010100001101000101",
"01000101010011100010110101000101",
"11111111110101001100011001010111",
"00101001000110100001101010000010",
"00001000000000000001101001000010",
"00000010010110101000010001000110",
"11111111010001100001110100001110",
"10000100010001100001110000001111",
"10000000010001100000000101011010",
"01010110000101100000111100001010",
"00110101010000000000000100001111",
"01011010100000000100011000000000",
"00010110000011110000111100000010",
"00101101010000000000000001000110",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"01011010100000000100011000001000",
"00011010100000000100011000000001",
"00001111000010100001011000001111",
"00001001100100001001000101010110",
"01010110000000000000100001000000",
"00011010000110100001000000001111",
"10101101100110000000000100010110",
"11110010110000101001111110111000",
"11000110000010101000100111111111",
"00111101100000011111111111010100",
"01011000010001010000000000001110",
"01010100010101010100001101000101",
"01000101010011010010110101000101",
"01000100010011110100100001010100",
"10000010111111111101010011000110",
"00010111000110101000000001000110",
"01000010001010100010110101001110",
"00001010100100010000000000000100",
"01000110000010001000100000010000",
"00111000001011010100000000000000",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"00000001010110101000000001000110",
"10000001111111111101010011000110",
"01010110000000000000100100111101",
"01001111010011000100110001000001",
"01000101010101000100000101000011",
"10000010111111111101010011000110",
"00000000000001000100001000101011",
"00011010100000000100011000001000"
)
,(
"10001000010001100011011000001111",
"00011100001101100000001001011010",
"00001111000000000000110101000010",
"00010111010101010000001000001110",
"00000000000000110100001000101100",
"00001000000000010000111101010100",
"11111111110101001100011000000001",
"00000000000001110011110110000001",
"01010110010101000100010101010011",
"11000110010100000100111101010100",
"01010110100000101111111111010100",
"00000001000010100110000001000110",
"01011010100010000100011001010111",
"01011010100000000100011000000001",
"11010100010001100101010100000010",
"10000000010001100000000111111111",
"10000000010001100001011000011010",
"01000010010111000010110100001010",
"00000010000011100000000000011100",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"01000000000111010000100010000001",
"01010110000010011111111111011111",
"10010000000000100100000100111110",
"00010001000010011000001010010001",
"10010001010101101000100100010000",
"00000010000011100000100110010000",
"01000010001011000001011101010100",
"00001000100100000000000100000101",
"00000010000111010001000000011000",
"00000010000101100101011000001110",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"01010010000011100000100010000001",
"00001111001101010000001000010110",
"00101100000101110101010100000010",
"00000000000010110100001000011100",
"10000010111111111101010011000110",
"11000110000000010000111101010100",
"00001000100000011111111111010100",
"00000010000101100100111000001110",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"11000110100100000000100010000001",
"10000010100101100000000000010100",
"11111111111111111000110110001110",
"11000010100111000000000000000000",
"01000110000011100000000001100101",
"00000010000101100000000000100000",
"00000000001010000100011000001111",
"00001111001101010000001000010110",
"00110110000101110101001000000010",
"00000000010010110100001000011100",
"10000010111111111101010011000110",
"11000110000000010000111101010010",
"00010000100000011111111111010100",
"00000000111111111111111100001101",
"00111000000110010001110000000000",
"00000000000100000100011000010000",
"00111000000101110101000000100011",
"00000000001010110100001000100010",
"01010110000011110000001000011101",
"01000000000010011001000010010001",
"00000010000011100000000000011010",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"10011000000111010000100010000001",
"11000010100111111011100010101101",
"00001001100010011111111111100000",
"01000110000000000010111001000000",
"00001110000101100000000000011000",
"10010000100100010101011000000010",
"00000000000110100100000000001001",
"00110101000000100000111000011101",
"00010111010101010000001000001111",
"00001011010000100001110000101100",
"11111111110101001100011000000000",
"00000001000011110101010010000010",
"10000001111111111101010011000110",
"10111000101011011001100000001000",
"11111111111000001100001010011111",
"10001001000100010000100010001001",
"10000010111111111101010011000110",
"11000110000000010000111101010010",
"00011101100000011111111111010100",
"10111000101011011001100000011101",
"11111110111010101100001010011111",
"01000010001011000000100010001001",
"00010111001111101111111011010101",
"01010110000000100000111100000001",
"00001110000010011001000010010001",
"00101100000101110101010100000010",
"00001110000000000000010101000010",
"00001000000001000110000100111110",
"10101101100110000001110100011101",
"11101010110000101001111110111000",
"01000110000010011000100111111111",
"00001000000000101111111111010100",
"01011010100010000100011001010110",
"00000000111011000011111000000001",
"10010001010101100000001000001111",
"00000010000011100000100110010000",
"00001010001101100010110101001110",
"00001010000111000011011000001111",
"01010101000000000000001101000010",
"00011101000111010000000100001111",
"10011111101110001010110110011000",
"10001001111111111110011111000010",
"11111111110101001100011000001001",
"00000000000000100011110110000001",
"11011100001111100010000101010110",
"11011000001111101001000000000000",
"11111111111111000000110100000101",
"01010101000000100000010111111111",
"10001000000100000010000000010000",
"00011010000110100001011101010011",
"11011101001111100001011000011010",
"00001010010110000100011000000101",
"10001000000100000000000110010000",
"00110001001111100000000100011101",
"00111110010100100011110100000000",
"00000010000010011111011001110011",
"00111101111111111100111100111110",
"01010010010000110000000000001000",
"01000101010101000100000101000101",
"01011000010001100100110101001101",
"01000010001101010000001000001010",
"00001101000011100000000000000111",
"00000101111111111111111111111100",
"00001110000101110000111000000001",
"10010000000010100101100001000110",
"00011101100010000001000000000001",
"01011000010001100011110100000001",
"00000010000111011001000000001010",
"00110101000000101000100000010000",
"00001111000000000011010101000010",
"00000001000111010001110100001111",
"00010000010101010000111010010001",
"00010000000011100001011000100000",
"00011010000101110101001110001000",
"00001111000000000101000100111110",
"00001111000011110000000100001111",
"01010110000010000000000100011101",
"00001111010101100000000100001111",
"00001111010011000000000100011101",
"00011101000000100001010000111110",
"00000000111111100100011000011101",
"01010110000000000011010100111110",
"00000001000010100110000001000110",
"00000000000010010011110100001001",
"01000101010011000100010101010010",
"01001101010001010101001101000001",
"10010000100100010101011001001101",
"00000000000010110100000000001001",
"00000001000011110000001000001111",
"00011101000010001001000000011101",
"10101101100110001000100000010000",
"11101111110000101001111110111000",
"00111101000010011000100111111111",
"00000010000010100101100001000110",
"00111101000111010001110100001110",
"00001001100100001001000101010110",
"01010110000000000000010101000000",
"10011000000111010000000100001111",
"11000010100111111011100010101101",
"00001000100010011111111111110101",
"00000000000111111100011000111101",
"00111000000100000001111100101001",
"00000000000001010100001000011100",
"11110011010000000001101010011001",
"00011000001011000001101011111111",
"00111101000101101000100000010000",
"00001010001010100010110101010001",
"00001000000000000000001001000010",
"00001010010110001100011000111101",
"10010000100000101001110100010000",
"00001110000110011000001000001000",
"00011010001000010001011100010001",
"01010101000100000001101000011010",
"00010110000101100010000000010001",
"00000010000111010000111010010001",
"01010101000101110001000100001110",
"00101100001001000010000000010000",
"00001000000000000001000001000010",
"00010001000011100000001000001110",
"00100000000100000101010100010111",
"00000010010000100010110000100100",
"00001111010101100000100000000000",
"00010000000000100001110110010000",
"00110110000101110000001010001000",
"01000010000111000011011000001111",
"00001110100100010000000000101100",
"10101111001111101000100000010000",
"00010111000100010000111000000010",
"00100100001000000001000001010101",
"00010000010101010001011000010001",
"00011010001111100000111100100000",
"00010111000100010000100000000000",
"00011111001000000001000001010101",
"00001111000101100001000100011100",
"00010111000110100001101001010100",
"01010101001111100001100000010000",
"00001000000010010000111000000010",
"10010001001111011000100110001000",
"00001010010110001100011010010000",
"10010000100000101001110100010000",
"01000010000011111000001000001000",
"11010100010001100000000001000011",
"00001110000010000000001011111111",
"00111000001011010101001100000010",
"00100000010001100000111100001010",
"00011100001010100001011100000000",
"00000000000110110100001000101100",
"00011101000111010000111000001000",
"00010001010101010001000000000010",
"00010001000011110001011000100000",
"00011010000110100010000100010111",
"00001010100100010001011000011010",
"00000010010010000011111010010001",
"01010101100010010001000100010000",
"00000001111111111101010001000110",
"00001001100100001101010110010001",
"00010111100101100001000010100000",
"10111001010000001000100000010000",
"00010001100010010000100111111111",
"01000010000011111000100100010000",
"11010100010001100000000001011111",
"00001110000010000000001011111111",
"00111000001011010101001100000010",
"00100000010001100000111100001010",
"00011100001010100001011100000000",
"10010000000000000011001101000010",
"00000010000111010000111110010001",
"00000000100001010011111000001111",
"00000000000100100100001000110101",
"10101010001111100000111100010001",
"01000010001101010000101000000000",
"00011101100100000000000000001000",
"00000001000111010000111100011101",
"00110101000010101000100000010000",
"00010000000000000000101001000010",
"01010100000100010101010100001111",
"10010100001111100010000000010111",
"01000000100010010000100011111110",
"00001110000010000000000000000101",
"01010101000000100001110100011101",
"00000001111111111101010001000110",
"00001001100100001101010110010001",
"00010111100101100001000010100000",
"10011101010000001000100000010000",
"11010100010001100000100111111111",
"00111101000010000000001011111111",
"10000010000010100101100011000110",
"10001111110101010001000010001110",
"00001110100101101010000010000010",
"00010000000011110011011000000010",
"01000010000111000010101000010111",
"00011010010101000000000000000111",
"11101110010000000001011000011010",
"00010111000100000000111011111111",
"00000000000101110100001000101100",
"10010000000000100001000101010101",
"00010010001111100000111100100000",
"00010000010101010000111011111111",
"00111110001000000001011101010100",
"10001000000100001111111001011110",
"10001001000000010001000100011000",
"00001010010110001100011000111101",
"10010000100000101001110100010000",
"01010101000100001000001000001000",
"00001111000101100010000000010001",
"10010000001000010001011100010001",
"00010110000110100001101000011010",
"00000010000011110011011000010000",
"00001000010000100001110000101100",
"00011010000110100101010000000000",
"11101111010000001001100100010111",
"00001010000000100001110111111111",
"10010000001111011000100110001000",
"11000110100000101001110110011101",
"10011101000100000000101001011000",
"10000010000010001001000010000010",
"00100000000100010101010100001111",
"10001010000100010001011000010000",
"00011010000110100001011100010001",
"00001010100100010001011000011010",
"00110111001111100000111100001111",
"00010001100010100001000100000001",
"00001001100100001001000110001010",
"10010001000100011000100000010000",
"00010110010000100011011000010111",
"00011010000110100101010000000000",
"00010001000011111001100100010110",
"00100000000100000101010100010111",
"00001111000101100001000100100100",
"00000000110111100011111000010000",
"00001000111111111110000101000000",
"10001001000100000000000110010000",
"00001000100100000011110110001001",
"11111111011111010011111000001110",
"00000000000010000100001000101011",
"11111011001111110011111000001000",
"11111111011100010011111000001110",
"00000000000010010100001000101011",
"11101011001111100000111000001000",
"01100100001111100000111011111101",
"00001100010000100011010111111111",
"11111111100010110011111000000000",
"00000100010000100011010100001110",
"00011101000011110001000000000000",
"00111101000010101000100000000001",
"00101011000000000001100100111110",
"00001111000000000000010101000010",
"00001000000000010000111101001110",
"01000010000000000000110100111101",
"01000110010101000101001101000101",
"01000010010001010100010101010010",
"01001011010000110100111101001100",
"00000000010100000100001000110101",
"10000010111111111101010011000110",
"00011100010110100001011001001011",
"00001010011000000100011000001110",
"01100000010001100001011000000010",
"10001000001111100000000100001010",
"11111110110111000011111011111101",
"00000000000100110100001000110101",
"10001101001111100000111100001111",
"00001001010000100011010111111111",
"00001111000111010001110100000000",
"00001111010101010000000100011101",
"10010001000010100000111000000001",
"00110110100010000001000000001010",
"01000010000111000011011000001111",
"00011101000011100000000000010010",
"01010100000011110101010100000010",
"00000010000101110001101000011010",
"01010100001000000001011101010100",
"11111101001111000011111000010111",
"10000001111111111101010011000110",
"00000000000010000011110100101011",
"01001111010011000100110001000001",
"01000101010101000100000101000011",
"00000010000010100101100001000110",
"10011100110011111001000000010111",
"00011011000110110001101110101100",
"00011001100111001011100010010000",
"00001010010111000100011001010101",
"00100000000101110101001100000010",
"10001000000100000010101000010111",
"00000000000001100011110100011100",
"01001100010011000100000101001101",
"00001000100100000100001101001111",
"10011101100100001000001010010000",
"00011101000011110000111110000010",
"01000010001011000001000100000001",
"00001111000011110000000000000011",
"00001111000100000000100000000001",
"00001111010101100000000100011101",
"00000011010000100001000000000001",
"00000001000100000000111000000000",
"10011101000010001001000010001001",
"00001011001111011000000110011101",
"01001110010000010100100000000000",
"01010110010001010100110001000100",
"01000100010010010100110001000001",
"10011101100100011000001010010001",
"00000110010000100001000010000010",
"00000001000100000001000100000000",
"00010001000000000000001101000000",
"01000010000100010000000100001111",
"00010001000100000000000000000111",
"00000100010000000000000100011101",
"00011101000011110001000000000000",
"00111101000010011000100100000001",
"10000010111111111101010011000110",
"11111111011110000011111000001110",
"00110110000000100001110100001111",
"01101011010000100000111000011100",
"01010110000011100000111100000000",
"11000110110101100000000100001111",
"10011101000100000000101001011000",
"10000010000010001001000010000010",
"10010000000111010000111011010110",
"10000001000101110100111000000010",
"00100000000100010101010100010000",
"00010001000000100000111100010110",
"00011010001000010001011110010001",
"00001111000101100001101000011010",
"00010000010101010001011100010001",
"00010110000100010010010000100000",
"00101101010100110000001000001110",
"01000110000011110000101000111000",
"00101010000101110000000000100000",
"00001111001011000000101000011100",
"00010000000000100001110100011101",
"01000010000111000010110000010111",
"00111110000011110000000000011001",
"00010001000011111111111101111110",
"00100000000100000101010100010111",
"00010110000100010001110000011111",
"00010000000010100000101010010001",
"10011000000101110100111010001000",
"00001000111111111100010001000000",
"00101101001111101000100000010000",
"10001000000100001000100111111111",
"11111111110101001100011000001010",
"00111110000011110011110110000001",
"10001110010000101111111011111010",
"11111111110101001100011000000000",
"01011010000101100101001110000010",
"00000010000111010000111100011100",
"00010111000110100001101001010100",
"00100000000011110101010100000010",
"00001111000010100001011101001110",
"00000100010000100011100000101101",
"00010000000010101001000100000000",
"11111000001111100000100010001000",
"00101101000111000101101000000000",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"10010000000110110001101100001000",
"00000010000111010000111100001000",
"11111111111111111111110000001101",
"00010110010100110000001000000101",
"00111110000100000001110001011010",
"10000010100100011111101110111011",
"00000001000011110101010100001111",
"00001000111111110010100100111110",
"11100100001111100001011001001110",
"00001111000011110000111111111011",
"00110101111111011110111100111110",
"00011101000000000000100101000010",
"00000001000111010000111100011101",
"00001110000000010000111100010000",
"00001010100100011000100000001010",
"00001111001101101000100000010000",
"00010001010000100001110000110110",
"11111111111111000000110100000000",
"01010011000000100000010111111111",
"00001111000111000101101000010110",
"00111110000100000000001000011101",
"00101100100010001111101101111011",
"10000001111111111101010011000110",
"00001010000000000000010001000000",
"00111101111111011110100100111110",
"01010010010001100000000000000100",
"11010100110001100100010101000101",
"00111110000011101000001011111111",
"00010100010000101111111001010110",
"01010100000000100001110100000000",
"00000010000101110001101000011010",
"00010000000010101001000101010101",
"00011010010101000010000010001000",
"00000010010000000001011100011010",
"11000110000101110000111000000000",
"00111101100000011111111111010100",
"01000101010100100000000000000110",
"01000101010110100100100101010011",
"10000010111111111101010011000110",
"11111110001010000011111000001110",
"00001110000000000000010101000010",
"00000001000011110001100000000010",
"11111111110101001100011000001000",
"00000000000011100011110110000001",
"01001111010011000100110001000001",
"01000101010101000100000101000011",
"01001001010100110010110101000100",
"11010100110001100100010101011010",
"00111110000011101000001011111111",
"00010000010000101111111000000010",
"01010101000000100000111000000000",
"00100101010101101001000000010111",
"11000010101011000000000100001111",
"01101111001111100000000000000011",
"11010100110001100000100011111110",
"00001100001111011000000111111111",
"01000011010011100100100100000000",
"01000101010001100100010101010010",
"01000011010011100100010101010010",
"11111111110110000000110101000101",
"00001101000000100000010111111111",
"00000101111111111111111111111100",
"00001100001111010001011100000010",
"01000011010001010100010000000000",
"01000101010001100100010101010010",
"01000011010011100100010101010010",
"11111111111111000000110101000101",
"01010011000000100000010111111111",
"00001101000111000101101000010110",
"00000101111111111111111111111100",
"00000000000001100011110100000001",
"01010011010101010100111001010101",
"11111100000011010100010001000101",
"00000010000001011111111111111111",
"11111111111111000000110100010110",
"00111101000000010000010111111111",
"01001100010000010000000000000101",
"01000111010011100100011101001001",
"01000110110011110101100100111110",
"10001111001111100000000000010101"
)
,(
"11111111101010010011111011001111",
"01010101111100010010010100111110",
"00000010000010100101110001000110",
"00111110000110100010000000011001",
"00000000000011011111000100011010",
"00001101000010000000000000000000",
"00000101111111111111111111001100",
"00001011001111100001011100000010",
"00000000000110100100011011110001",
"00111101110011110010110100111110",
"01001100010000010000000000000101",
"01010000010101000100111101001100",
"00111101000111000101001100111101",
"01010010010101000000000000010000",
"01000101010001110100011101001001",
"01011001010100110010110101010010",
"01001111010011000100001101010011",
"00111101010100100100101101000011",
"01010010010101000000000000010001",
"01000101010001110100011101001001",
"01010010010100000010110101010010",
"01000001010000110101001101000101",
"01001111010100100100010101001100",
"01010100000000000000110100111101",
"01000111010001110100100101010010",
"01001001001011010101001001000101",
"01010100010101010101000001001110",
"00010110010011000001110001010011",
"10101011001111100000111100001111",
"00100000000011110101010111001101",
"00000010111111111101000001000110",
"11111111110100000100011000100010",
"00001100001111010000100100000001",
"01000011010011110100110000000000",
"01001111010000110010110101001011",
"01000101010101000100111001010101",
"00011010000110100001101001010010",
"00011010000110100000111100100010",
"00010110111111111100000001000110",
"00010011001111010000100000000001",
"01010100010001010101001100000000",
"01010101010011110100001100101101",
"01010010010001010101010001001110",
"01010010010001010101001100101101",
"01000101010000110100100101010110",
"11000000010001100001101000011010",
"00111101000000100001011011111111",
"01000101010100110000000000001010",
"01010101010011110100001101010100",
"01010010010001010101010001001110",
"00000010111111111101010001000110",
"00010000000010100110010011000110",
"00010000000000100001110110010000",
"01010101010101100000001010001000",
"00010000000101100000101010010001",
"00010000001001010000101010010001",
"10010000100010000001000010001001",
"00011101100010000001000000000001",
"11011000010001100000111000000001",
"11010100010001100000000111111111",
"01011100010001100000000111111111",
"00100000010001100000001000001010",
"00001010010110110010110100000000",
"01010101000000000000010001000010",
"01010100000010100010000000001111",
"00001010011000000100011000100011",
"01000110010110110001011100000010",
"00101100000000100101101010001000",
"00000000000000110100001000011100",
"00111101111101110001000000111110",
"01000101010100100000000000001011",
"01001111010000110100010001000001",
"01000101010101000100111001010101",
"01010011000000000000100001010010",
"01001100010000110101001101011001",
"00001001010010110100001101001111",
"01010101010011110101001100000000",
"00101101010001010100001101010010",
"00000000000001000100010001001001",
"01100010011010010111010000100011",
"01101001001111100000000000000011",
"01110100000000000000001101101110",
"00000000000000110110001001101001",
"00000011010001000100110001001000",
"01000100010000010101000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000"
)
                           );
  type dvec is array (0 to 9 - 1) of DataVec;
  signal bdata: dvec;
  signal old: std_ulogic_vector(ROMrange'high downto 11);
  
begin
  
  fetch: process(Clock) is
  begin
    if rising_edge(Clock) then
         old <= Address(old'range);
	   for i in bdata'range loop
	     bData(i) <= ROM(i)(to_integer(std_ulogic_vector(Address(11 - 1 downto 2))) MOD blocks'length);
		end loop;
	 end if;
  end process fetch;

  Data <= 
          bdata(0 ) when unsigned(old) = 0 else
          bdata(1 ) when unsigned(old) = 1 else
          bdata(2 ) when unsigned(old) = 2 else
          bdata(3 ) when unsigned(old) = 3 else
          bdata(4 ) when unsigned(old) = 4 else
          bdata(5 ) when unsigned(old) = 5 else
          bdata(6 ) when unsigned(old) = 6 else
          bdata(7 ) when unsigned(old) = 7 else
          bdata(8 ) when unsigned(old) = 8 else
          (others => '0');
			 
end RTL;
