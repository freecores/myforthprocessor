----------------------------------------------------------------------------------
-- Company: RIIC
-- Engineer: Gerhard Hohner Mat.nr.: 7555111
-- 
-- Create Date:    01/07/2004 
-- Design Name:    Diplomarbeit
-- Module Name:    ROMcode - Rtl 
-- Project Name:   32 bit FORTH processor
-- Target Devices: Spartan 3
-- Tool versions:  ISE 8.2
-- Description: implements a ROM containing the BIOS
-- Dependencies: global.vhd
-- 
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------


library IEEE, work;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.global.all;

entity ROMcode is
  port (Clock: in std_ulogic;									-- system clock
        Address: in std_ulogic_vector(ROMrange);		-- address bus
		  Data: out DataVec);									-- outgoing data
end ROMcode;

architecture RTL of ROMcode is
  type blocks is array (0 to 2048 / 4 - 1) of DataVec;
  type myarray is array (natural range <>) of blocks;
  constant ROM: myarray := (
(
"01000110010011100101011001010100",
"11100101001111100010010110000000",
"00000000000110110100011000100111",
"00000001111111111111000001000110",
"00111001000000000001011101000110",
"00000000000110000100011000000001",
"00001110010101100000000100110100",
"10010000000010100110110001000110",
"00011101100010000001000000000001",
"00111011001111100101001100000001",
"01000110000000100101101001000011",
"01100001001111100000001111101000",
"01000011100111110011111000010010",
"00000010111111111101010001000110",
"00101000000101110011111000001000",
"00001101001001111010111100111110",
"00000011000000000000000000000000",
"11111111111111111101100000001101",
"01000110010101100000000100000010",
"01010110000000010000101001000000",
"00000001000010100100010001000110",
"01100000010001100000111001010110",
"00010000000000011001000000001010",
"01010110000000010001110110001000",
"00000001000010101000000001000110",
"00001010100001000100011001010110",
"10011000010001100101011000000001",
"01000110010101100000000100001010",
"01010110000000010000101010010000",
"00000001000010101001010001000110",
"00001010100010000100011001010110",
"10001100010001100101011000000001",
"01000110010101100000000100001010",
"01000110000000010000101001101000",
"00001101010100100000101010101100",
"00000100000000000000110100111110",
"00000000000011000101100100111110",
"01010010010101100000000000000000",
"00000000000011010011100000001101",
"00001100010011000011111000000100",
"01001100000000000000000000000000",
"00001101001100100000110101010010",
"00111111001111100000010000000000",
"00000000000000000000000000001100",
"00000000000000000000000000001101",
"00101001000011010101001000000011",
"00111110000001000000000000001101",
"00000000000000000000110000101110",
"00000000000000000000110100000000",
"00001101010100100000001100000000",
"00000100000000000000110100011110",
"00000000000011000001110100111110",
"00010000010001100000000000000000",
"00010011000011010101001000000000",
"00111110000001000000000000001101",
"00000000000000000000110000001110",
"00001010011011000100011000000000",
"00001101000001010000110101010010",
"11111111001111100000010000000000",
"00000000000000000000000000001011",
"00000000000011001110110000001101",
"01110101000011010101001100000100",
"00111110000001000000000000001101",
"11000001000011010000101111101110",
"01010011000001000000000000001101",
"00000000000011100001001000001101",
"00001011111000000011111000000100",
"00000000000011011100110100001101",
"01110110000011010101001100000100",
"00111110000001000000000000001110",
"00011000000011010000101111010010",
"01010011000001000000000000001110",
"00000000000011101100011100001101",
"00001011110001000011111000000100",
"00000000000011101101000000001101",
"11011100000011010101001100000100",
"00111110000001000000000000001110",
"11010110000011010000101110110110",
"01010011000001000000000000001110",
"00000000000011101110101100001101",
"00001011101010000011111000000100",
"00000000000011101110011100001101",
"00011111000011010101001100000100",
"00111110000001000000000000001111",
"11110110000011010000101110011010",
"01010011000001000000000000001110",
"00000000000011110010100100001101",
"00001011100011000011111000000100",
"00000000000011110010010100001101",
"10100010000011010101001100000100",
"00111110000001000000000000001111",
"11110000000011010000101101111110",
"01010011000001000000000000001111",
"00000000000100000011110000001101",
"00001011011100000011111000000100",
"00000000000100000111000000001101",
"10011100000011010101001100000100",
"00111110000001000000000000010000",
"10000110000011010000101101100010",
"01010011000001000000000000010000",
"00000000000100001100101000001101",
"00001011010101000011111000000100",
"00000000000100001010001000001101",
"11010101000011010101001100000100",
"00111110000001000000000000010000",
"11010000000011010000101101000110",
"01010011000001000000000000010000",
"00000000000100001111100000001101",
"00001011001110000011111000000100",
"00000000000100001101110100001101",
"00010011000011010101001100000100",
"00111110000001000000000000010001",
"11111111000011010000101100101010",
"01010011000001000000000000010000",
"00000000000100011011110000001101",
"00001011000111000011111000000100",
"00000000000100010001011100001101",
"11010011000011010101001100000100",
"00111110000001000000000000010001",
"11000011000011010000101100001110",
"01010011000001000000000000010001",
"00000000000100011110000100001101",
"00001011000000000011111000000100",
"00000000000100011101110000001101",
"00001111000011010101001100000100",
"00111110000001000000000000010010",
"11101001000011010000101011110010",
"01010011000001000000000000010001",
"00000000000100100010110100001101",
"00001010111001000011111000000100",
"00000000000100100001011100001101",
"01110010000011010101001100000100",
"00111110000001000000000000010010",
"00110101000011010000101011010110",
"01010011000001000000000000010010",
"00000000000100100111111100001101",
"00001010110010000011111000000100",
"00000000000100100111101000001101",
"10001111000011010101001100000100",
"00111110000001000000000000010010",
"10000011000011010000101010111010",
"01010011000001000000000000010010",
"00000000000100101001011100001101",
"00001010101011000011111000000100",
"00000000000100101001001000001101",
"10100010000011010101001100000100",
"00111110000001000000000000010010",
"10011101000011010000101010011110",
"01010011000001000000000000010010",
"00000000000100101011000000001101",
"00001010100100000011111000000100",
"00000000000100101010010100001101",
"10111010000011010101001100000100",
"00111110000001000000000000010010",
"10110101000011010000101010000010",
"01010011000001000000000000010010",
"00000000000100111000111100001101",
"00001010011101000011111000000100",
"00000000000100101100000100001101",
"10100011000011010101001100000100",
"00111110000001000000000000010011",
"10010011000011010000101001100110",
"01010011000001000000000000010011",
"00000000000100111111111100001101",
"00001010010110000011111000000100",
"00000000000100111010110000001101",
"01001111000011010101001100000100",
"00111110000001000000000000010100",
"00001000000011010000101001001010",
"01010011000001000000000000010100",
"00000000000101001001110100001101",
"00001010001111000011111000000100",
"00000000000101000101011100001101",
"00011111000011010101001100000100",
"00111110000001000000000000010101",
"10100101000011010000101000101110",
"01010011000001000000000000010100",
"00000000000101010110010000001101",
"00001010001000000011111000000100",
"00000000000101010010011100001101",
"10100000000011010101001100000100",
"00111110000001000000000000010101",
"01101000000011010000101000010010",
"01010011000001000000000000010101",
"00000000000101011010111100001101",
"00001010000001000011111000000100",
"00000000000101011010010000001101",
"11111001000011010101001100000100",
"00111110000001000000000000010101",
"10110101000011010000100111110110",
"01010011000001000000000000010101",
"00000000000101100101001000001101",
"00001001111010000011111000000100",
"00000000000101100101011100001101",
"00100101000011010101001100000100",
"00111110000001000000000000010111",
"00101101000011010000100111011010",
"01010011000001000000000000010111",
"00000000000110000011101100001101",
"00001001110011000011111000000100",
"00000000000110000111000000001101",
"01100100000011010101001100000100",
"00111110000001000000000000011001",
"01011101000011010000100110111110",
"01010011000001000000000000011001",
"00000000000110110000111100001101",
"00001001101100000011111000000100",
"00000000000110010110100000001101",
"01111010000011010101001100000100",
"00111110000001000000000000011011",
"00010011000011010000100110100010",
"01010011000001000000000000011011",
"00000000000111000000001100001101",
"00001001100101000011111000000100",
"00000000000110110111111000001101",
"01010001000011010101001100000100",
"00111110000001000000000000011100",
"00001111000011010000100110000110",
"01010011000001000000000000011100",
"00000000000111000111111000001101",
"00001001011110000011111000000100",
"00000000000111000101011000001101",
"10100110000011010101001100000100",
"00111110000001000000000000011100",
"10000110000011010000100101101010",
"01010011000001000000000000011100",
"00000000000111001100110000001101",
"00001001010111000011111000000100",
"00000000000111001010110100001101",
"11111011000011010101001100000100",
"00111110000001000000000000011100",
"11010010000011010000100101001110",
"01010011000001000000000000011100",
"00000000000111010001000100001101",
"00001001010000000011111000000100",
"00000000000111010000000100001101",
"00101101000011010101001100000100",
"00111110000001000000000000011101",
"00011001000011010000100100110010",
"01010011000001000000000000011101",
"00000000000111010100110000001101",
"00001001001001000011111000000100",
"00000000000111010011001000001101",
"01100100000011010101001100000100",
"00111110000001000000000000011101",
"01010011000011010000100100010110",
"01010011000001000000000000011101",
"00000000000111011000100100001101",
"00001001000010000011111000000100",
"00000000000111010110110000001101",
"10101010000011010101001100000100",
"00111110000001000000000000011101",
"10010000000011010000100011111010",
"01010011000001000000000000011101",
"00000000000111011111101100001101",
"00001000111011000011111000000100",
"00000000000111011011000100001101",
"00101011000011010101001100000100",
"00111110000001000000000000011110",
"00000011000011010000100011011110",
"01010011000001000000000000011110",
"00000000000111100101100100001101",
"00001000110100000011111000000100",
"00000000000111100011001000001101",
"10101100000011010101001100000100",
"00111110000001000000000000011110",
"01100001000011010000100011000010",
"01010011000001000000000000011110",
"00000000000111101101001000001101",
"00001000101101000011111000000100",
"00000000000111101011010000001101",
"00011011000011010101001100000100",
"00111110000001000000000000011111",
"11011000000011010000100010100110",
"01010011000001000000000000011110",
"00000000000111110010111100001101",
"00001000100110000011111000000100",
"00000000000111110010001000001101",
"11010000000011010101001100000100",
"00111110000001000000000000011111",
"00110101000011010000100010001010",
"01010011000001000000000000011111",
"00000000000111111110010100001101",
"00001000011111000011111000000100",
"00000000000111111101100000001101",
"11111011000011010101001100000100",
"00111110000001000000000000011111",
"11101010000011010000100001101110",
"01010011000001000000000000011111",
"00000000001000000100110000001101",
"00001000011000000011111000000100",
"00000000001000000000001000001101",
"01110000000011010101001100000100",
"00111110000001000000000000100000",
"01010010000011010000100001010010",
"01010011000001000000000000100000",
"00000000001000001000001000001101",
"00001000010001000011111000000100",
"00000000001000000111011000001101",
"11011100000011010101001100000100",
"00111110000001000000000000100000",
"10001001000011010000100000110110",
"01010011000001000000000000100000",
"00000000001000001110110000001101",
"00001000001010000011111000000100",
"00000000001000001110010100001101",
"00010101000011010101001100000100",
"00111110000001000000000000100001",
"11110011000011010000100000011010",
"01010011000001000000000000100000",
"00000000001000010100001100001101",
"00001000000011000011111000000100",
"00000000001000010001101100001101",
"10101010000011010101001100000100",
"00111110000001000000000000100001",
"01001010000011010000011111111110",
"01010011000001000000000000100001",
"00000000001000011011010100001101",
"00000111111100000011111000000100",
"00000000001000011010111000001101",
"11011100000011010101001100000100",
"00111110000001000000000000100001",
"10111010000011010000011111100010",
"01010011000001000000000000100001",
"00000000001000011110011100001101",
"00000111110101000011111000000100",
"00000000001000011110000000001101",
"00011101000011010101001100000100",
"00111110000001000000000000100010",
"11101101000011010000011111000110",
"01010011000001000000000000100001",
"00000000001000100010100100001101",
"00000111101110000011111000000100",
"00000000001000100010001000001101",
"01001110000011010101001100000100",
"00111110000001000000000000100010",
"00101111000011010000011110101010",
"01010011000001000000000000100010",
"00000000001000100110011000001101",
"00000111100111000011111000000100",
"00000000001001001100100100001101",
"11100001000011010101001100000100",
"00111110000001000000000000100100",
"11010101000011010000011110001110",
"01010011000001000000000000100100",
"00000000001001001111000000001101",
"00000111100000000011111000000100",
"00000000001001001110010100001101",
"00011100000011010101001100000100",
"00111110000001000000000000100101",
"11110110000011010000011101110010",
"01010011000001000000000000100100",
"00000000001001010010110100001101",
"00000111011001000011111000000100",
"00000000001001010010001000001101",
"00111111000011010101001100000100",
"00111110000001000000000000100101",
"00110000000011010000011101010110",
"01010011000001000000000000100101",
"00000000001001010110111000001101",
"00000111010010000011111000000100",
"00000000001001010111001000001101",
"10000100000011010101001100000100",
"00111110000001000000000000100101",
"01111101000011010000011100111010",
"01010011000001000000000000100101",
"00000000001001011000111100001101",
"00000111001011000011111000000100",
"00000000001001011000101000001101",
"10101011000011010101001100000100",
"00111110000001000000000000100101",
"10010100000011010000011100011110",
"01010011000001000000000000100101",
"00000000001001011011011000001101",
"00000111000100000011111000000100",
"00000000001001011010111100001101",
"11000000000011010101001100000100",
"00111110000001000000000000100101",
"10111011000011010000011100000010",
"01010011000001000000000000100101",
"00000000001001011100100100001101",
"00000110111101000011111000000100",
"00000000001001011100010000001101",
"11101001000011010101001100000100",
"00111110000001000000000000100101",
"11001100000011010000011011100110",
"01010011000001000000000000100101",
"00000000001001011111010000001101",
"00000110110110000011111000000100",
"00000000001001011110110100001101",
"00000100000011010101001100000100",
"00111110000001000000000000100110",
"11111010000011010000011011001010",
"01010011000001000000000000100101",
"00000000001001100001010000001101",
"00000110101111000011111000000100",
"00000000001001111110111000001101",
"10101101000011010101001100000100",
"00111110000001000000000000101000",
"01010011000011010000011010101110",
"01010011000001000000000000101000",
"00000000001010001110000000001101",
"00000110101000000011111000000100",
"00000000001010001110100000001101",
"10000011000011010101001100000100",
"00111110000001000000000000101001",
"00010011000011010000011010010010",
"01010011000001000000000000101001",
"00000000001010011100001000001101",
"00000110100001000011111000000100",
"00000000001010011000100100001101",
"11010110000011010101001100000100",
"00111110000001000000000000101001",
"11000111000011010000011001110110",
"01010011000001000000000000101001",
"00000000001010011110111000001101",
"00000110011010000011111000000100",
"00000000001010011101110000001101",
"00000111000011010101001100000100",
"00111110000001000000000000101010",
"11110101000011010000011001011010",
"01010011000001000000000000101001",
"00000000001010100001110100001101",
"00000110010011000011111000000100",
"00000000001010100001011000001101",
"00110000000011010101001100000100",
"00111110000001000000000000101010",
"00101001000011010000011000111110",
"01010011000001000000000000101010",
"00000000001010100111100100001101",
"00000110001100000011111000000100",
"00000000001010100011011100001101",
"10010011000011010101001100000100",
"00111110000001000000000000101010",
"10000001000011010000011000100010",
"01010011000001000000000000101010",
"00000000001010101111000100001101",
"00000110000101000011111000000100",
"00000000001011101110111000001101",
"11110011000011010101001100000100",
"00111110000001000000000000101110",
"11110000000011010000011000000110",
"01010011000001000000000000101110",
"00000000001011101111101000001101",
"00000101111110000011111000000100",
"00000000001011101111100000001101",
"00000001000011010101001100000100",
"00111110000001000000000000101111",
"11111111000011010000010111101010",
"01010011000001000000000000101110",
"00000000001011110000100000001101",
"00000101110111000011111000000100",
"00000000001011110000011000001101",
"00101101000011010101001100000100",
"00111110000001000000000000101111",
"00001101000011010000010111001110",
"01010011000001000000000000101111",
"00000000001011110100011000001101",
"00000101110000000011111000000100",
"00000000001011111011001000001101",
"00111011000011010101001100000100",
"00111110000001000000000000110000",
"01000111000011010000010110110010",
"01010011000001000000000000110000",
"00000000001100000101010100001101",
"00000101101001000011111000000100",
"00000000001100000101000000001101",
"10001100000011010101001100000100",
"00111110000001000000000000110000",
"01100010000011010000010110010110",
"01010011000001000000000000110000",
"00000000001100001110011100001101",
"00000101100010000011111000000100",
"00000000001100001001011100001101",
"01000100000011010101001100000100",
"00111110000001000000000000110001",
"11110100000011010000010101111010",
"01010011000001000000000000110000",
"00000000001100010101010100001101",
"00000101011011000011111000000100",
"00000000001100010101001100001101",
"10001010000011010101001100000100",
"00111110000001000000000000110001",
"01100000000011010000010101011110",
"01010011000001000000000000110001",
"00000000001100011011010000001101",
"00000101010100000011111000000100",
"00000000001100011011111000001101",
"00000110000011010101001100000100",
"00111110000001000000000000110010",
"11001000000011010000010101000010",
"01010011000001000000000000110001",
"00000000001100100110011000001101",
"00000101001101000011111000000100",
"00000000001100100111000100001101",
"11011110000011010101001100000100",
"00111110000001000000000000110010",
"11110000000011010000010100100110",
"01010011000001000000000000110010",
"00000000001100110100101000001101",
"00000101000110000011111000000100",
"00000000001100110001110100001101",
"10001010000011010101001100000100",
"00111110000001000000000000110011",
"01011011000011010000010100001010",
"01010011000001000000000000110011",
"00000000001100111011111000001101",
"00000100111111000011111000000100",
"00000000001100111001011100001101",
"11111011000011010101001100000100",
"00111110000001000000000000110011",
"11001100000011010000010011101110"
)
,(
"01010011000001000000000000110011",
"00000000001101000101001000001101",
"00000100111000000011111000000100",
"00000000001101000000011100001101",
"10101111000011010101001100000100",
"00111110000001000000000000110100",
"01011110000011010000010011010010",
"01010011000001000000000000110100",
"00000000001101001011111100001101",
"00000100110001000011111000000100",
"00000000001101001011110000001101",
"00010100000011010101001100000100",
"00111110000001000000000000110101",
"11001101000011010000010010110110",
"01010011000001000000000000110100",
"00000000001101010110010000001101",
"00000100101010000011111000000100",
"00000000001101010111000100001101",
"01111111000011010101001100000100",
"00111110000001000000000000110101",
"01111000000011010000010010011010",
"01010011000001000000000000110101",
"00000000001101011110111100001101",
"00000100100011000011111000000100",
"00000000001101011000111000001101",
"00011001000011010101001100000100",
"00111110000001000000000000110110",
"11111101000011010000010001111110",
"01010011000001000000000000110101",
"00000000001101100100101100001101",
"00000100011100000011111000000100",
"00000000001101100010100100001101",
"01110010000011010101001100000100",
"00111110000001000000000000110110",
"01010001000011010000010001100010",
"01010011000001000000000000110110",
"00000000001101101001111100001101",
"00000100010101000011111000000100",
"00000000001101100111100100001101",
"11010100000011010101001100000100",
"00111110000001000000000000110110",
"10101110000011010000010001000110",
"01010011000001000000000000110110",
"00000000001101110000111000001101",
"00000100001110000011111000000100",
"00000000001101101110000000001101",
"01000100000011010101001100000100",
"00111110000001000000000000110111",
"00011010000011010000010000101010",
"01010011000001000000000000110111",
"00000000001101111000000100001101",
"00000100000111000011111000000100",
"00000000001101111000100100001101",
"00111011000011010101001100000100",
"00111110000001000000000000111000",
"10110000000011010000010000001110",
"01010011000001000000000000110111",
"00000000001110011010010000001101",
"00000100000000000011111000000100",
"00000000001110000100101000001101",
"00000011000011010101001100000100",
"00111110000001000000000000111010",
"10110001000011010000001111110010",
"01010011000001000000000000111001",
"00000000001110100110011100001101",
"00000011111001000011111000000100",
"00000000001110100001001100001101",
"10011010000011010101001100000100",
"00111110000001000000000000111010",
"01110010000011010000001111010110",
"01010011000001000000000000111010",
"00000000001110101100110100001101",
"00000011110010000011111000000100",
"00000000001110101010010100001101",
"11000101000011010101001100000100",
"00111110000001000000000000111100",
"11010110000011010000001110111010",
"01010011000001000000000000111010",
"00000000001111001111100100001101",
"00000011101011000011111000000100",
"00000000001111001100100100001101",
"00001111000011010101001100000100",
"00111110000001000000000000111101",
"00011001000011010000001110011110",
"01010011000001000000000000111101",
"00000000001111011000000100001101",
"00000011100100000011111000000100",
"00000000001111011100010000001101",
"01110111000011010101001100000100",
"00111110000001000000000000111110",
"11111001000011010000001110000010",
"01010011000001000000000000111111",
"00000000010000000011101000001101",
"00000011011101000011111000000100",
"00000000010000000010101100001101",
"10011111000011010101001100000100",
"00111110000001000000000001000000",
"01001001000011010000001101100110",
"01010011000001000000000001000000",
"00000000010000001100111100001101",
"00000011010110000011111000000100",
"00000000010000001010100100001101",
"00000000000011010101001100000100",
"00111110000001000000000001000001",
"00110001000011010000001101001010",
"01010011000001000000000001000001",
"00000000010000100101100100001101",
"00000011001111000011111000000100",
"00000000010000011011001000001101",
"10000101000011010101001100000100",
"00111110000001000000000001000010",
"01011111000011010000001100101110",
"01010011000001000000000001000010",
"00000000010000101010001100001101",
"00000011001000000011111000000100",
"00000000010000101000110100001101",
"11010100000011010101001100000100",
"00111110000001000000000001000010",
"10110011000011010000001100010010",
"01010011000001000000000001000010",
"00000000010000101111000000001101",
"00000011000001000011111000000100",
"00000000010000101110001000001101",
"00001111000011010101001100000100",
"00111110000001000000000001000011",
"11111110000011010000001011110110",
"01010011000001000000000001000010",
"00000000010000110010010100001101",
"00000010111010000011111000000100",
"00000000010000110001011100001101",
"01011101000011010101001100000100",
"00111110000001000000000001000011",
"01100100000011010000001011011010",
"01010011000001000000000001000011",
"00000000010000110110100100001101",
"00000010110011000011111000000100",
"00000000010000110110011000001101",
"01111101000011010101001100000100",
"00111110000001000000000001000011",
"01111011000011010000001010111110",
"01010011000001000000000001000011",
"00000000010000111001001000001101",
"00000010101100000011111000000100",
"00000000010000111001000000001101",
"11000101000011010101001100000100",
"00111110000001000000000001000011",
"10100001000011010000001010100010",
"01010011000001000000000001000011",
"00000000010000111110000100001101",
"00000010100101000011111000000100",
"00000000010000111101001100001101",
"11111110000011010101001100000100",
"00111110000001000000000001000011",
"11110110000011010000001010000110",
"01010011000001000000000001000011",
"00000000010001000111011100001101",
"00000010011110000011111000000100",
"00000000001111001111100100001101",
"00000000001111100101011000000100",
"00001010010101000100011000000011",
"01000100110010110000110100000001",
"00111110010101100000010000000000",
"01011000010001100000001011110011",
"01000000010001100000000100001010",
"11000110000011010101010100001000",
"00111110000001000000000001000100",
"10101000010001100000001001010010",
"11000001000011010101010100001010",
"00111110000001000000000001000100",
"01000000010001100000001001000110",
"10111100000011010101010100001001",
"00111110000001000000000001000100",
"01001000010001100000001000111010",
"10110111000011010101010100001001",
"00111110000001000000000001000100",
"01001100010001100000001000101110",
"10110001000011010101010100001001",
"00111110000001000000000001000100",
"01010101010101100000001000100010",
"00000000010001001010011000001101",
"00000010000110000011111000000100",
"00001101010101010000001001011010",
"00000100000000000100010010011100",
"01000110000000100000110100111110",
"00001101010101010000101001011000",
"00000100000000000100010011001011",
"01000110000000100000000100111110",
"00001101010101010000101001010100",
"00000100000000000100010010010101",
"01000110000000011111010100111110",
"00001101010100100000101010010000",
"00000100000000000100010010001100",
"01000110000000011110100100111110",
"00001101010100100000101010001100",
"00000100000000000100010010000100",
"01000110000000011101110100111110",
"00001000000000101111111111010100",
"00000000000000000000110101010110",
"00010100000000000000010000000000",
"01000110001100100001111000111110",
"00001000000000101111111111010100",
"11110000000000001000110111010110",
"10010100100000000000001111111111",
"01000110000001000100000001000110",
"01000110000000010000100101000000",
"01000100010001100000010000000000",
"01000110010101100000000100001001",
"01010110000000010000101010011100",
"00000001000010101010000001000110",
"00001010101001000100011001010110",
"01001100010001100101011000000001",
"01000110010101010000000100001010",
"01010110000000010000101001010000",
"00000001000010010100100001000110",
"00001001010011000100011001010110",
"01011100010001100101011000000001",
"00000000010001100000000100001010",
"00001001010001000100011000000100",
"00000100010000000100011000000001",
"00000001000010010100000001000110",
"11111111110100000100011001010111",
"00000000000100000100011000000001",
"00001001100100001001000101010110",
"11111111110110000100011000001110",
"10111000101011011001100000000001",
"11111111111101001100001010011111",
"00100110000110110000110110001001",
"00111110010010010000010000000000",
"00001001000011010000001100111110",
"01001000000001000000000000100110",
"00001101000000110011010100111110",
"00000100000000000100010000001010",
"00000011001011000011111001000111",
"00000000000011110011000000001101",
"00100011001111100101011000000100",
"11111111110100000100011000000011",
"00011111111111100100011000000010",
"11111111110100000100011000011100",
"00011110010110100011111000000001",
"00001010010010000100011001010110",
"11010100010001100101010100000001",
"00011111001111100000000111111111",
"11000010000011010000100000011101",
"00011110000001000000000000001110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"10010011001111100010001000000100",
"00101100001111100101010100000100",
"11111111110101000100011000100011",
"01001000010001100000100000000010",
"01000110010101100000001000001010",
"01010101000000010000101001001000",
"00000001111111111101010001000110",
"00100011000101010011111001010111",
"00000000111111110100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"11011100010000001111010000101110",
"11111110010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000110001000010",
"00001010100000000100011001010110",
"00100001011001110011111000000001",
"00000000000000001100011001000000",
"00101101000000001111110101000110",
"00000111010000100000101000101100",
"01100001001111100000100000000000",
"00000000101101010100000000101001",
"00000000111111000100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000001000",
"01000000000010000001110010101010",
"01000110000000000000000010100011",
"00101100001011010000000011111011",
"00000000000001110100001000001010",
"00000010101001100011111000001000",
"00000000000000001001001001000000",
"00101101000000001111101001000110",
"00000111010000100000101000101100",
"01010100001111100000100000000000",
"00000000100000010100000000011100",
"00000000111110010100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"01110000010000000011011010111010",
"11111000010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000011101000010",
"01000000001100001000001000111110",
"01000110000000000000000001011111",
"00101100001011010000000011110111",
"00000000000001110100001000001010",
"00110000100001010011111000001000",
"00000000000000000100111001000000",
"00101101000000001111011001000110",
"00000111010000100000101000101100",
"10011000001111100000100000000000",
"00000000001111010100000000110000",
"00000000111101010100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"00101100010000000000000111001000",
"11110100010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000011101000010",
"01000000001000010111010100111110",
"01000110000000000000000000011011",
"00101100001011010000000011110011",
"00000000000100000100001000001010",
"00000000000000000000110100001000",
"10000000010001101000000000000000",
"10100010001111100000000100001010",
"00000000000000010100000000100000",
"11111110111101010100000000001000",
"00000000000000000000000000111101",
"11111111111111111101100010001101",
"11010011100000101000111000000010",
"10001110100101111001101010011010",
"00010000100111010000000100010000",
"10001000000100001001110100000001",
"10001000100000011000111100000001",
"01001101000000000000110000111101",
"01001001010011000100110001001001",
"01001111010000110100010101010011",
"00001001010100110100010001001110",
"01000101010100100101000000000000",
"01001001010100110100100101000011",
"00000000000010010100111001001111",
"01010101010001000100111101001101",
"01001111010101000100010101001100",
"01000100000000000000011101010000",
"01010100010101000100001101001001",
"00000000000001000101000001001111",
"01000101010100110100000101000010",
"01010000010100110000000000000100",
"00000000000001000100111001000001",
"01000101010100100100010101001000",
"00011001000011100001111000001110",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"10010001010101100001111000001010",
"00000100000011110000100110010000",
"00110101000101110000010000001111",
"00001010000000000000010001000010",
"00001000001111011000100100001010",
"00011000000010001001000000011000",
"10101101100110001000100000010000",
"11100101110000101001111110111000",
"01010110000010011000100111111111",
"01100011000000000000011000111101",
"01110100011000010110010101110010",
"00000000000000000000110101100101",
"11011000000011010000001100000000",
"00000010000000101111111111111111",
"01000000000010011001000010010001",
"00010001100100000000000000101000",
"11111111010001100000001000011101",
"00101101000100000001110000000000",
"10001000000100000000101000101100",
"01000010000111000010001000101100",
"00010000000011110000000000001110",
"11111111100111000011111000000010",
"00000000000001000100001000101100",
"00111101100010010001000000001001",
"10010000000110100001101001010011",
"10111000101011011001011000001000",
"11111111110100101100001010011111",
"00010111000011100000100010001001",
"00111110010101100000111000111101",
"01000010001101011111111110110111",
"00110101000010100000000000000010",
"11111111111100010011111000111101",
"01010110000000000000010001000010",
"00001000000000010001110100001111",
"00000000000000000000010000001101",
"00000000000000000000110100000011",
"11011000000011010000001100000000",
"00000010000000101111111111111111",
"00001001100100001001000100011101",
"00010000000000000001000101000000",
"00000000000001100100001000000010",
"01000000100010010001000000001000",
"00011010010100110000000000001101",
"10010110000010001001000000011010",
"11000010100111111011100010101101",
"01010101100010011111111111101001",
"00001101000101110001101000011010",
"00000010111111111111111111011000",
"00000000000001000011110100000001",
"01000100010011100100100101000110",
"10010000000111010000111100110110",
"00000000111111110100011000000010",
"10000010100111010001110000011100",
"00101100001011010101011000000000",
"00000000000001110100001000001010",
"00111101100010000000100000001000",
"00000000000000000011111101000000",
"00001010001011000010110101010011",
"00001000000000000000011001000010",
"00110001010000000011110100001000",
"00101101010100010000000000000000",
"00010100010000100000101000101100",
"11001100100011010000100000000000",
"10000001000000101111111111111111",
"00001101000111010001110100011101",
"00000010111111111111111111011000",
"00010101010000000011110100000001",
"00101101010100000000000000000000",
"00001100010000100000101000101100",
"11111100100011010000100000000000",
"10000001000000101111111111111111",
"00000001010000000011110100001000",
"00010000000010000000100000000000",
"00000000000001100011110110001000",
"01100111011100100110111101100110",
"00111110010101110111010001100101",
"00101100000010100010001110001011",
"00000000000010110100001010010000",
"11110000001111100101000100001110",
"10011100100100000011010111111110",
"00001000111111111000010100111110",
"11000010000000100100011000111110",
"11000010000011010000000000001000",
"01000000000001000000000000001110",
"10111001000011010000000000000101",
"00111110000001000000000000001110",
"00001110000111100000001000110011",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000001101110000011111000100010",
"01000110000000000000011100111101",
"01000101010011000100100101000001",
"00000000000000110011111001000100",
"00000111001111100100101101001111",
"01000101010110000100010100000000",
"01000101010101000101010101000011",
"00011010000110100001110001000111",
"00011100010001110011110100000001",
"00111101000000100001101000011010",
"01000101010100110000000000001001",
"01000011010001010101011001010100",
"00111110010100100100111101010100",
"00001001001111011111110000110101",
"01010100010001010100011100000000",
"01010100010000110100010101010110",
"01001111010001100101001001001111",
"00011110010000100000010000001010",
"11111001001111100100011100000000",
"00000000000101000100011000000000",
"01010110000000010011110000111110",
"01000110001000111011010100111110",
"11101001001111100000000000011001",
"00001010011101000100011000000000",
"11111111111111000000110100000010",
"00111110000000010000001011111111",
"00000100001111011111101111110001",
"01001001010101010101000100000000",
"00000001000011100101101001010100",
"01000001000000000000010100111101",
"01010100010100100100111101000010",
"11111111110101000100011001000011",
"00001111011111010000110100000010",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000001001010000011111000100010",
"11111111111111111110010000001101",
"00010000010001100000001000000010",
"11111111111001000000110100000000",
"00010000000000010000001011111111",
"00001101000101100010111100111110",
"00000010111111111111111111100100",
"11011000010001100000111000000001",
"11010100010001100000000111111111",
"01000000000011010000000111111111",
"01010110000000000000111101000010",
"10011000000010011001000010010001",
"11000010100111111011100010101101",
"01000100100010011111111111111001",
"01110101000000000010001100111101",
"01100110011001010110010001101110",
"01100100011001010110111001101001",
"01110011011011100110100100100000",
"01100011011101010111001001110100",
"01101110011011110110100101110100",
"01100011011011110110110000100000",
"01100100011001010111010001100001",
"01100001011001010110111000100000",
"00000000000001110010000001110010",
"01010100010001100100111101010011",
"01000110010101000100111001001001",
"11000110000000101111111111010100",
"01000100110001100000101001000000",
"00010000000000100001000100001010",
"00000000000110000100011000000010",
"00000010111111111110110001000110",
"00101100000101110001110000001111",
"01000010000111000011100000001111",
"00010111010101000000000000011100",
"00000000010000000100011000001111",
"11100000010001100000011000010110",
"00001010100100010000000111111111",
"01000110000111101000100000010000",
"10010001000111000000001111111111",
"01000000100010000001000000001010",
"00000001000100001111111111010011",
"01000110100010010000000100010001",
"00111101000000011111111111010100",
"00000010000010100100010001000110",
"00010111000001000000000001000110",
"11110011001111100011110100101010",
"11111111111110100100001011111111"
)
,(
"01000110000000000001100001000110",
"00001111000000101111111111101100",
"01000110001011000001011100011100",
"00101100000000100000101001000100",
"00000000000001110100001000011100",
"00000001111111111110000001000110",
"11000110000000000010000001000000",
"11000110100000101111111111010100",
"10000010100011100000101001000100",
"00000010000010100100000001000110",
"11111111010001100001011000010000",
"01000000010001100001110000000011",
"10011110000001010001011000000000",
"11000110100010001000000110001111",
"00111101100000011111111111010100",
"01001101010001010000000000000101",
"01000110001111110101010001001001",
"00001110000111000000000011111111",
"00010111000000000001101101000110",
"00000100010000100001111100111000",
"00000001000000000100011000000000",
"11111111101000100011111000100010",
"10010000100100010101011000111101",
"00000000000001110100000000001001",
"11011110001111100000010000001110",
"10101101100110000001100011111111",
"11110011110000101001111110111000",
"00111101000010001000100111111111",
"00011110100110010011111001010101",
"11111111100000100011111001010110",
"01000110111111111101111000111110",
"01111001001111100000000000011010",
"10001000001111100101011111111111",
"00111110010101010011110100011110",
"00111110010101100001111010000011",
"10110010001111101111111101101100",
"00000000000110100100011011111111",
"01010111111111110110001100111110",
"00111101000111100111001000111110",
"01011001010101000000000000000100",
"00111110010101010100010101010000",
"00111110010101100001111001100111",
"10010001010101101111111101010000",
"00000111010000000000100110010000",
"00000000001000000100011000000000",
"10011000111111111000110000111110",
"11000010100111111011100010101101",
"01000110100010011111111111110011",
"00110101001111100000000000011010",
"01000100001111100101011111111111",
"00000000000001000011110100011110",
"01010100010010010100110101000101",
"11111111110011100011111001010101",
"01010011000000000000011000111101",
"01000101010000110100000101010000",
"00101100001111100101010101010011",
"00010101001111100101011000011110",
"01011010001111100100100111111111",
"01010110001111100100110011111111",
"00000000000110100100011011111111",
"01010111111111110000011100111110",
"00111101000111100001011000111110",
"01010000010100110000000000000101",
"01010101010001010100001101000001",
"01010110000111100000101000111110",
"00111110001001010100101000111110",
"00111110010101111111111101100110",
"00111110010101110010010101000011",
"00000010001111010001110111111011",
"00001111010100100100001100000000",
"01000010001011000010001000001111",
"00001010000010000000000000001000",
"00011001000011100000111000001010",
"10011000110101100011110100001110",
"00001111000010011001000010010001",
"10010001000100000001000100001111",
"10010001000100000001011100001010",
"10001001000100000010011000001010",
"01000011000100000001000100001001",
"00101010100010010001000100011111",
"00001010010000100001110000011111",
"10011010000010001001000000000000",
"10001000000100000010010100001110",
"00010000111111111101100001000000",
"00110101100011101101011010001000",
"00011001000000000010011001000010",
"10010000100100010000100010010000",
"00010000000101110000101010010001",
"00010000001001100000101010010001",
"01000010000111110100001110001001",
"01010101000100010000000000110110",
"00101000010101010001000000100011",
"10001001000100010001000010001001",
"00011000101001011000111000011010",
"11010110010000000000100010010000",
"01000000000010010000100011111111",
"01000010001101010000000000110110",
"10010000000110010000000000101000",
"00100011010101010000100110010001",
"00101000010101011000100000010000",
"00001010100100011001000010010001",
"00001010100100010001000000010110",
"01000011100010010001000000100101",
"11111111110010100100001000011111",
"00010000100010010001000000010001",
"10001110000110101000100100010001",
"01000000000010001001000010100101",
"10010001000010001111111111010100",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00111101100010010001000000010001",
"01010010010100000000000000000101",
"10010000010101000100111001001001",
"10001000000100000001011100001110",
"10010001111111110100110000111110",
"00010001000010100000100110010000",
"00000111001111011000100100010000",
"00101111010001000101010100000000",
"01000100010011110100110101000100",
"00001010111111111110010000111110",
"01010101000000000000011000111101",
"01001111010011010010111101000100",
"10010001000010001001000001000100",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"00101001000100011000100000010000",
"00100001000000000000000101000010",
"10100100111111111101100100111110",
"00000000000001101100001010101010",
"00100001000010001001000000100001",
"00000110001111011000100000010000",
"00101111010011010101010100000000",
"10010000010001000100111101001101",
"10010000111111111100111000111110",
"00001001010000100010100100001000",
"01000010001010100001000100000000",
"00010001001000010000000000000001",
"10001001000100001001100100010110",
"01010011000000000000011000111101",
"01000101010100100010111101001101",
"00001001100100001001000101001101",
"01000010001010010001000001010110",
"00010001001000010000000000000001",
"00000000000000010100001000101001",
"00100000010001101010010000100001",
"10010000100100010101011000000000",
"00011011100100001001000100001001",
"00010110000111000010011000001110",
"00010000000100010010100001010101",
"10011000100010010010100001010101",
"11000010100111111011100010101101",
"00001010100010011111111111101011",
"00000000000010011100001010101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00000000000001100011110110001000",
"01001101001011110100110101000110",
"10111000001111100100010001001111",
"00000010001111010000101011111111",
"10010000001010100100110100000000",
"00010000001010101001000000001000",
"00111110100010000001000010001000",
"00000001001111011111111101011011",
"11101110001111100010101000000000",
"00000100001111010000101011111111",
"01001111010011010010111100000000",
"11111111111000110011111001000100",
"00000000000000010011110100001000",
"00111110000010001001000000101111",
"10001000000100001111111110001011",
"00111101111111110011101000111110",
"01001111010011010000000000000011",
"11111111111011010011111001000100",
"00000000000001010011110100001010",
"01001111010011010010111100101010",
"01000110000001000000111101000100",
"00101100001011010000000000101101",
"00000000000001010100001000001010",
"00000111010000001000111011010111",
"11000110100100001101011000000000",
"10101100100101110000000000101011",
"00000000000001101100001000001000",
"00011000000010001001000000011001",
"00001000100100001000100000010000",
"00000000100100111100001010110111",
"00110000010001100000010010010000",
"00001010001010100010110100000000",
"00000000001110010100011000001111",
"00011111001000100011100000010111",
"00011100000000000011000001000110",
"00000000010000010100011000010111",
"00001111000010100010101000101101",
"00010111000000000101101001000110",
"01000110000111110010001000111000",
"00010111000111000000000000110111",
"00101101000000000110000101000110",
"01000110000011110000101000101010",
"00111000000101110000000001111010",
"01010111010001100001111100100010",
"00001101000101110001110000000000",
"00000010111111111111111111100100",
"00011111001010100010110100000010",
"00001001000000000000011001000010",
"01000110010000001000100000010000",
"00001001100100001001000100000000",
"01010110000010011001000010010001",
"10001001000100000001000100001110",
"00000000001000111100001010110101",
"00100110000011100000111010011011",
"10010001000000000000111001000010",
"00010110000010101001000110010000",
"00100101000010101001000100010000",
"00010000000100011000100100010000",
"10010001000011110000111110001001",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00001001111111111101100101000000",
"10010001100010010001000100010000",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"10011001000110001000100000010000",
"00010001111111110110100101000000",
"01000010000010101001000110001010",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"00010000100010000001000000001010",
"00000010001111011000100100010001",
"00011110001011110010101000000000",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"00100000001111100010001000000100",
"00000111001111010000100011111111",
"01010101010011100011111000000000",
"01010010010001010100001001001101",
"00000000000001110100001000101001",
"00000000010101000011111000100001",
"01000110000000000100011101000000",
"00111000001011010000000001000000",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"10101010100100010000100010010000",
"00011111010001101000101000010001",
"01000010001110000010110100000000",
"00011001000101110000000000001110",
"10010001000100010000100110010000",
"00010000100010000001000000001010",
"11111111111010100100000010001000",
"00001111001000111001000000001000",
"00010000000000000010000001000110",
"10010001001000100010000000010111",
"00010000100010000001000000001010",
"00100000010001100001000100100011",
"00010111100010010001000000000000",
"00001010100100010010001000100000",
"00000111001111011000100000010000",
"01001110010011110100001100000000",
"01010100010100100100010101010110",
"00000000000001110100001000101001",
"11111111100111000011111000100001",
"01000110000000000011101101000000",
"00111000001011010000000001000000",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"00101101000000000001111101000110",
"00000000000011110100001000111000",
"00001000100100000001100100010111",
"10001000000100000000101010010001",
"10001000000100000001011100001110",
"00001000111111111110100101000000",
"10010001001000001001000110010000",
"00010001100010000001000000001010",
"00100000010001100001000000100000",
"00100011000101110001000100000000",
"00010000000010101001000100100010",
"00000110001111011000100110001000",
"01001000010100110100000100000000",
"00101001010101000100011001001001",
"00100001000000000000011101000010",
"01000000111111111010100100111110",
"01000000010001100000000000111010",
"01000010001110000010110100000000",
"00001010100100010000000000000100",
"01000110000010001000100000010000",
"00111000001011010000000000011111",
"00010111000000000000111101000010",
"00001110000010001001000000011001",
"00010000000010101001000100010111",
"01000000100010000001000010001000",
"10010000000010001111111111101001",
"00100000010001100000111100100011",
"00100000000101110001000000000000",
"00010000000010101001000100100010",
"00100011100010000001000010001000",
"10001000000100000000101010010001",
"01010011000000000000011000111101",
"01010100010001100100100101001000",
"00101010000011111001000101001100",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"10010001000010011001000010010001",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10001010000100011000100000010000",
"10010001100100001000101000010001",
"00001001100100011001000000001001",
"01000000010001100000111001010110",
"00110100010000100011010100000000",
"00001000100100000001100100000000",
"00001110000010001001000000011010",
"00010001100010000001000000100101",
"10001001000100000001000110001010",
"10001110100010000001000010011010",
"10010001000010001001000010100101",
"00010001100100010000100010010000",
"01000011000010001001000010001010",
"10010001000000000000110001000010",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00001001000000000000000101000000",
"11001000010000001000100000010000",
"10001001100010010000100011111111",
"00001001110000101010101010100100",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"00000110001111011000100000010000",
"01001001010010000101001100000000",
"10010001010100100101010001000110",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10010001100100001000100000010000",
"00101010000011111001000100001001",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"10001010000100011000101000010001",
"11111011110001110011111010100100",
"00000000000010011100001010101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00001010000010001001000010001000",
"00111101100010000001000000001010",
"00101010010001000000000000000010",
"01000010001010100000111110010001",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"10010000100010000001000000001010",
"00001111100100010000100110010001",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00010001100010100001000110001000",
"10000110001111101010010010001010",
"11000010101010100000100111111011",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"00111101100010000001000000001010",
"00101111010001000000000000000010",
"00000000000011010000100010010000",
"00100100100000000000000000000000",
"00000100001111011000100000010000",
"01001111010011010100010000000000",
"00100010000011110000111101000100",
"00000000000000010100001000101100",
"01000010001010100000111100111101",
"00111111110001100000000000001111",
"00001000100100000010000100001100",
"00001010001001100000111101010110",
"00000011010000001000100000010000",
"00000100001111111100011000000000",
"10010001000011110000111110011001",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"11111111111100000100001001000011",
"01000110000011110010001101001010",
"00100010001000000000000000010100",
"00100011010010100000100010010000",
"00000000000101000100011000010001",
"10001001000100000010001000100000",
"01000110000000000000011100111101",
"01000001010001110100010101001110",
"00001000100100000100010101010100",
"00001101000010011001000010010001",
"00111111111100000000000000000000",
"00010000100010111101010001010110",
"00000001010000100010100110001000",
"01000010000011100010000100000000",
"01000011000110110000000000100010",
"00010001000000000000100101000010",
"00111110000100010000101010010001",
"10001000000100000000000100000111",
"00001010100100011000101000010001",
"00001111000011111000101000010001",
"10010001000000001111101000111110",
"10010001100010100001000100001010",
"11111111110110100100000000001010",
"11000010101010101000100100001000",
"10010000100100010000000000001111",
"00000000000000000000110100001001",
"00010001010101100011111111110000",
"00010111001111101000100100010000",
"00000000000000110011110100000011",
"10010000010001100011111001000100",
"00001110010101100000100110010001",
"00111110100010010001000100010000",
"00001111100100001111110001011111",
"00000000001011100100011000000100",
"00110110000011110010110000010111",
"00000000001100100100001000011100",
"00001000100100000001100110001000",
"10010001000010001001000000011000",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10001010000100011000100000010000",
"11111100001101010011111000010001",
"10001010000100010000100010010000",
"01000010001010100000101010010001",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"00010000100010000001000000001010",
"10010111100100001000100100010001",
"00001001100100011001000010100001",
"00010000111111110000101000111110",
"00000000010001010100011000000100",
"00001111000010100010110000101101",
"00010111000000000110010101000110",
"00010001000010100010001000101100",
"00010000010000100001110000110110",
"00010000000011100101011000000000",
"10001001000110010001000100011000",
"00001001111110111111011000111110",
"10010001100100001001011010010000",
"00001101010101101000100100001001",
"00000010111111111111111111100100",
"11111110110110010011111000000010",
"00100001001111101000100000010000",
"00000000010010010011111011111111",
"00110101010001100011110101010111",
"10010000100100010101011000000000",
"10010000100110111001000100001001",
"10010000000010011010100011010101",
"10010000110000110000100110010001",
"10001000000100000001101100001000",
"00001000110000100010100001010101",
"10010000000101100001000100000000",
"00010000001001010001000100001000",
"10001001000100010001000010001000",
"10011000100010010001000000010001",
"11000010100111111011100010101101",
"00001001100010011111111111010111",
"00011011000010001001000000001001",
"10100101110101101010100011010101",
"10001000000100000010010101010110",
"00111110000000000000011000111101",
"01000001010011110100110001000110",
"10010000000010001001000001010100",
"00001111111111111111111110001101",
"00000000000011011001110000000000",
"00011100111111111111000000000000",
"00000000000000000000110100001110",
"00110110000111000111111111110000",
"10001101000000000000011001000010",
"00000000000100000000000000000000",
"10010001000010101001000110100010",
"11111111100011010001000000001010",
"10011100000000000000111111111111",
"11110000000000000000000000001101",
"00001101000011100001110011111111",
"01111111111100000000000000000000",
"00000110010000100011011000011100",
"00000000000000001000110100000000",
"10010000101000100000000000010000",
"00000000100011011010010010010001",
"10011100100000000000000000000000",
"11110000000000000000000000001101",
"10010001000110110001110001111111",
"00001101100010000001000000001010",
"01111111111100000000000000000000",
"00001101000101100001101100011100",
"00011111111110000000000000000000",
"00000000000000000000110100010111",
"00111000001011010011111111110000",
"00000000000011100100001000001010",
"00000000000011011001101000001000",
"01010101111111111110000000000000",
"10001001100010000101011000101000",
"00101101010101100011110110001001",
"00000000000001000100001000101010",
"10001000000100000000101010010001",
"00001000100100000001101000001000",
"00010001000011100101011010100010",
"00001111100010100001000110001010",
"00010110000010101001000100001111",
"00100101000010101001000100010000",
"10001010000100011000100100010000",
"00010101001111101000101000010001",
"00000000000011010000111111111111",
"00101101000000000001000000000000",
"00000110010000100000101000101010",
"00000000000000001000110100000000",
"00001101100111001000000000000000",
"00000000000111111111111111111111",
"00001101010000100011100000010111",
"00011011000010001001000000000000",
"10001000000100001010100011010101",
"00010000000000000000000010001101",
"00001000100100001001011000000000",
"00001111111111111111111100001101"
)
,(
"00100010000100010001110000000000",
"10010001001111011000100100010000",
"11111111000011010000100010010000",
"00011100000000000000111111111111",
"00000000000000000000110100010001",
"10010000000111000111111111110000",
"00001101000000000000011001000010",
"00000000000100000000000000000000",
"00011010100010100001000100100010",
"00100101000011100000100010010000",
"00101010000100011000100000010000",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00000010001111011000100100010000",
"01000110001010100100011000000000",
"00101010000101110000000000110010",
"00001010100100010000100010010000",
"00011010100010010001000000010001",
"00100011000000000001010101000110",
"00001010100100010000100010010000",
"00011010100010010001000000010001",
"00100011000000000001010101000110",
"00101001000101110000111100001111",
"00100001000000000000000101000010",
"00010111000000000011011001000110",
"00011100001101100000111100101010",
"00111101000111000000101000001010",
"00111110000010011001000010010001",
"10001010000100011111111110010001",
"10001010000100010000101010010001",
"10010000111111111000100000111110",
"00010100010001100001000100001000",
"01000110000100000010001100000000",
"00010111001000110000000000010100",
"00000000000011110100001000101001",
"10010001000010101001000110001010",
"00010011001111100010000100001010",
"10001001000100010001000011111011",
"10001000000000000000010001000000",
"10010001111110110000100100111110",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"11010101000110100000111110011010",
"00101010000011110000100010101000",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00101100001000100000111100001111",
"10001101000000000000011001000010",
"10000000000000000000000000000000",
"00000000000011010000111110011100",
"00010111000000000010000000000000",
"00011100000110100001000000101010",
"00001111000000000001010001000010",
"00010110000010101001000100001111",
"00100101000010101001000100010000",
"00000000100011011000100100010000",
"10010111000000000001000000000000",
"00010000111111111101111001000000",
"10010001010101100101010010001000",
"00001000100100000000100110010000",
"11111111111111110000110100001111",
"00111000000101110000000000111111",
"00000000000011010001101000010000",
"00010111111111111110000000000000",
"00001101010000100001110000110110",
"00011011000010001001000000000000",
"00101000010101011000100000010000",
"00010000000000000000000010001101",
"00001110010101101001011000000000",
"00010110000010101001000100011000",
"00100101000010101001000100010000",
"00011100010110001000100100010000",
"10101101100110001000100000010000",
"11000101110000101001111110111000",
"00001000100100001000100111111111",
"00010000000110110000100010010000",
"00001111001010000101010110001000",
"00001111111111111111111100001101",
"00010000001110000001011100000000",
"01000010000111000010110000011010",
"00000000100011010000000000000110",
"10010110000000000001000000000000",
"11111111000011010000100010010000",
"00011100000000000000111111111111",
"10001001000100000010001000010001",
"11111100010001000011111000111101",
"00111101111111110000110100111110",
"00101011010001100000000000000010",
"00100010000011110001101000001111",
"00000000000011100100001000101100",
"00011010001001000000101000001000",
"00000000000000000000110100001000",
"00101000010101011111111111100000",
"00001110000011110011110101010110",
"00001111111111111111111100001101",
"00001101000011110001110000000000",
"01111111111100000000000000000000",
"00000000000001100100001000011100",
"00010000000000000000000000001101",
"10010000000010100010001000000000",
"00001000100100000000100110010001",
"10001101100100011001000010010001",
"00000000000011111111111111111111",
"00000000100011011001000110011100",
"10011100011111111111000000000000",
"10001101000000000000011011000010",
"00000000000100000000000000000000",
"00001110010101100000100110100010",
"00010000100010010001000100010000",
"00000000000101010100011000011010",
"01000110000110100001000100100011",
"00010111001000110000000000010101",
"00010110000000111111111101000110",
"00000001000000000000000000001101",
"10001101101001000001011000000000",
"10000000000000000000000000000000",
"10100010000010001001000010011100",
"10001000000100000000111100001111",
"00010001000010101001000100010001",
"00010000000101110000101010010001",
"00010000001001100000101010010001",
"00011111001010100000100010001001",
"00010000000000000000110101000010",
"10001110000110101000100100010001",
"00001001100100011001000010100101",
"11111111110111000100000010011000",
"11111111111111110000110100010000",
"00001101000111000000000000000001",
"00000000000000010000011111111110",
"01000010000010100011100000101101",
"00001001000010010000000000001111",
"00000000000011011001101000001000",
"01010101111111111110000000000000",
"10001000100010010101011000101000",
"11111111110010110000110100111101",
"00101010001011010000000000000000",
"00000000000011100100001000001010",
"10001101000010000000100100001001",
"10000000000000000000000000000000",
"10001001010101100001000010011100",
"00000000000011010011110110001000",
"00101101000000000000000100000000",
"00001101010000100000101000101010",
"00000000000000001000110100000000",
"01000110100111001000000000000000",
"01000000001000100000000000000000",
"00010111000011100000000000000010",
"00010110000000000011011101000110",
"00000000000001111111111110001101",
"10001000000100001001110010000000",
"00001010100100011000101000010001",
"00001000100100001000101000010001",
"10001010000100010000101010010001",
"00000000001010011100001010110111",
"10010001100100001001000110011001",
"10010001000100000001011100001010",
"10001001000100000010011000001010",
"00101101010000100001111101000011",
"00001000100100000001101000000000",
"00001000100100000010010100001110",
"00001110000010001001000000011010",
"10001000000110000001000000100101",
"00010001100010010001000100010000",
"11010011010000001000100100010000",
"00101000110000101011011111111111",
"10010000100100011001100100000000",
"00010000000101100000101010010001",
"00010000001001010000101010010001",
"01000010000111110100001110001001",
"10010000000110101111111111010011",
"10010000001001010000111000001000",
"00001000100100000001101000001000",
"10001000000100000010010100001110",
"00010001100010010001000100010000",
"11010100010000001000100100010000",
"00001001000010011000100011111111",
"00001000100100001001000010010001",
"11010110101010001101010100011011",
"00010000001001010101011010100101",
"00000000000011010000111110001000",
"00011100000000000011000000000000",
"00010000000000000000000000001101",
"01000010001011000001011100000000",
"10011001100010010000000000000101",
"00001001000000000000111001000000",
"01010110100101101101010000010001",
"10101000110101010001101100100101",
"01010101100010010001000000011011",
"00001101000010001001000000101000",
"00000000000011111111111111111111",
"00010101010001100001000100011100",
"00011010000100010010000000000000",
"00100010001010000101010100001000",
"00000010001111011000100100010000",
"10010001001011010100011000000000",
"00010001010101100000100110010000",
"00000000000000000000000000001101",
"00011010000100010001110010000000",
"00100011000000000001010101000110",
"00010111000000111111111101000110",
"00000011111111100100011000011111",
"00000000000101010100011000010110",
"00100010001000110101010100100000",
"00001111010101101101011010010000",
"00111110000010110101001000010001",
"00011010000100011111110100000001",
"00100011000000000001010101000110",
"00010111000001111111111101000110",
"00100010010000100001110000101010",
"10001001000100000001000100000000",
"00001111111111010001110100111110",
"00001111000011110000111100001111",
"11111011110100010011111000001111",
"11001100001111100001000000010001",
"11111101111110010011111011111011",
"01010100000010011001000010010001",
"00001100010101000001100000001011",
"10010000111111111100100001000000",
"00010001000010101001000100001000",
"10001001000010001000100100010000",
"00000000000000100011110110001001",
"00001101000011110010111101000110",
"10000000000000000000000000000000",
"00000000000000000000110100011100",
"01010110001000100011111111100000",
"00111110111111001110000100111110",
"00000000000000000000000001111101",
"00000000000011010000111100000000",
"00011100011111111111000000000000",
"00100011000000000001010001000110",
"00010111000000111111111101000110",
"00000000000001110100001000101001",
"00001110010101100000100100001000",
"01000110000000000101001101000000",
"00111000001011010000000000111110",
"00000000000101110100001000001010",
"00001001010000100010101000001001",
"00000000000000000000110100000000",
"01000000010101101000000000000000",
"11111111000011010000000000000110",
"01010111011111111111111111111111",
"10010000000000000011001101000000",
"00001101100100000000100110010001",
"00000000000011111111111111111111",
"00000000000000000000110100011100",
"00010001001000100000000000010000",
"00110100010001100001000110001010",
"01000010001101110001011100000000",
"00011011001111100000000000000110",
"00000000000001000100000011111000",
"11111000011000110011111000100001",
"00000000000010011100001010101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00001010001111011000100010001000",
"01000011010001010101001000000000",
"01001111010100100101000001001001",
"00001111010011000100000101000011",
"11110000000000000000000000001101",
"00000000000011010001110001111111",
"00010111001111111111000000000000",
"00000000000010010100001000101001",
"00000000000000000000110100001001",
"01010110000111001000000000000000",
"00000000000101000100011000111101",
"00000000001101001100011000100011",
"10110111100101110000100010010000",
"01010111000000000001100011000010",
"10010111000000000010000011000110",
"00000000000010101100001010101001",
"00010000000000000010000001000110",
"01000000000111000010000000010110",
"00010000000010100000000000000101",
"10001000010101100001110000100000",
"01000110000000000000001100111101",
"00001111000011110100010000111110",
"10010001111111111011010000111110",
"10010001000010001001000010010000",
"00010000101001000010010000001010",
"00011111001011000010001010001000",
"00010001000111000010101000010001",
"00010001000010101001000110001010",
"00000000000010011100001010001010",
"11110000000000000000000000001101",
"11100000001111100101011000111111",
"00000000000001100011110111111100",
"01101001011100100111010001110011",
"00001111000011110110011001110000",
"00001011010100010000101101010001",
"00001111111111001100111000111110",
"00001111001101100010001000011010",
"00011111000010100001110000101010",
"10010001000000000000100101000010",
"00010001000010010000100110010000",
"00001111000011111000100100010000",
"00000000000001010011110100001001",
"01001111010011110100110001000110",
"01010001000011110000111101010010",
"00111110000010110101000100001011",
"00011010000011111111110010100111",
"00101010000011110011011000100010",
"00001001010000100000101000011100",
"00001001100100001001000100000000",
"10001001000100000001000100001001",
"00111101000010010000111100001111",
"01001101010001100000000000000100",
"00001111000011110101100001000001",
"10010001111111110011100000111110",
"10010001000010001001000010010000",
"00010000101001000010010000001010",
"00011111001011000010001010001000",
"00011100000111110010101000010001",
"00001010100100011000101000010001",
"00001001110000101000101000010001",
"00000000000000000000110100000000",
"00111110010101100011111111110000",
"00000100001111011111101101110110",
"01001001010011010100011000000000",
"00001001100100001001000101001110",
"00010001000000100010111000111110",
"00100000001111101000100100010000",
"00000001110010000011111011111010",
"01000110000000000000011000111101",
"01001110010101010100111101010010",
"00000000010100000011111001000100",
"11111001001000011111101100001101",
"00101101000110000000110100111111",
"00110100001111100101010001000100",
"11111000011110000011111011111100",
"01000110000000000000001100111101",
"00001111000011110010101000101010",
"11110100001111100000111100001111",
"00000000000000000000110111111001",
"00111110010101100011111111110000",
"01000100001111101111110000011011",
"11111011001010000011111000000011",
"00111101000000011110101000111110",
"01000001010001100000000000000101",
"00001101010100110100111101000011",
"01000000000000100110101110110001",
"10110101010101010001011100001101",
"11111001110011010011111010111011",
"00111101000000010111010100111110",
"01000001010001100000000000000110",
"01001000010100110100111101000011",
"00000000000011011001000010010001",
"01010110001111111111000000000000",
"00001111100010010001000000010001",
"11111001101100010011111000001111",
"00111110111110111101111000111110",
"11100011001111100000001100000111",
"00000000001010010011111011111011",
"01000110000000000000010100111101",
"01000111010011110100110001000001",
"00001111000011110000111100001111",
"00001101111110011001011000111110",
"00111111111100000000000000000000",
"11111010110100000011111001010110",
"00111110000000101110011000111110",
"10001100001111101111101011001010",
"00000000000001010011110100000001",
"01001001010100110100000101000110",
"00001111000011110000111101001110",
"11111001011101010011111000001111",
"10010001111101111110100100111110",
"10010000100100010000100110010000",
"00010000000100010101011000001001",
"00001011010100100001000100001111",
"01000010111110100111010000111110",
"00010000000100010000000000100010",
"00111110000100000001000110001001",
"10010000100100011111100101010111",
"00001110000110000000101101010010",
"00011000000110100000110001010001",
"10001000000100000010101010010000",
"00111110111101111100111000111110",
"10000011001111101111101101111110",
"11111111110101000100000011111010",
"00001010100100010000100010010000",
"00001000100010010001000000010001",
"00000110001111011000100110001001",
"01010011010000010100011000000000",
"01010011010010000100111001001001",
"10010001000010001001000000001011",
"00111110111110110101110100111110",
"11000010101010101111111110100011",
"11111011000011010000000000010111",
"00001101010000000000100100100001",
"01010100010001000010110100011000",
"00000000000001101100001010101001",
"01000000111110110011101000111110",
"01000111001111100000000000000011",
"00000101001111011000100011111010",
"01010100010000010100011000000000",
"00000000000011010100111001000001",
"01010110001111111111000000000000",
"00001111111110100011010100111110",
"00000000000000000000110100001111",
"00111110010101100100000000000000",
"01011011001111101111101100010111",
"11111011000111000011111011110111",
"00001101000000001110011000111110",
"00111111111000000000000000000000",
"11111000110101010011111001010110",
"01000110000000000000011000111101",
"01001110010000010101010001000001",
"00111110000011110000111100110010",
"00111011001111101111100011000111",
"00001001100100001001000111110111",
"00000000000000000000110101010110",
"10010001010101100011111111110000",
"01010010000100010000111110010000",
"11111001110000110011111000001011",
"00010001000000000010001001000010",
"00010000000100011000100100010000",
"01010010111110001010011000111110",
"01010001000011100001100000001011",
"00011001000011100001101000001100",
"00111110111100111010001000111110",
"11001111001111101111011100011111",
"00111110100100001001000111111010",
"11010100010000001111100111010010",
"10010001000010001001000011111111",
"10001001000100000001000100001010",
"00111101100010011000100100001000",
"01000001010001100000000000000110",
"01001000010011100100000101010100",
"10010001000000000010000100111110",
"00000000000000000000110110010000",
"00010001010101100011111111110000",
"10100011001111101000100100010000",
"11111001101010000011111011111010",
"11100000000000000000000000001101",
"01011100001111100101011000111111",
"00000000000001000011110111111000",
"01010011010011110100001101000110",
"10010000100100011001000010010001",
"00000000000011010101010100001001",
"01010110001111111111000000000000",
"10000111001111100001000000010001",
"01010010000100010000111111111001",
"11111001010011110011111000001011",
"00010001000000000001110101000010",
"00010000000100011000100100010000",
"01010110111110000011001000111110",
"00001110000110000000101101010001",
"10110000001111100000110001010000",
"11111010011000000011111011110110",
"01100011001111101001000010010001",
"11111111110110010100000011111001",
"00001010100100010000100010010000",
"00001000100010010001000000010001",
"00000101001111011000100110001001",
"01001111010000110100011000000000",
"10110011001111100100100001010011",
"00000000000000000000110111111111",
"00111110010101100011111111110000",
"00000100001111011111101000101111",
"01011000010001010100011000000000",
"00001101000011100000111101010000",
"01111111111100000000000000000000",
"00101010000011110010110000011100",
"00001100010000100000101000100010",
"00001000000110100000100000000000",
"11100000000000000000000000001101",
"01010110001010000101010111111111",
"00001000100100001001000100111101",
"00000000000101010100011000011010",
"00000011111111110100011000100011",
"00010000001010101001000000010111",
"11110110010100010011111010001000",
"11100110001011100100001000001101",
"00111001111011110000110100111111",
"10111100001111101111111011111010",
"00010001000100000001000111110111",
"00000000000000000000110110001001",
"01010110000111000111111111110000",
"10010001111110011110100100111110",
"00000000000000000000110110010000",
"00111110010101100011111111110000",
"00010000000100011111100111010011",
"11111001110110000011111010001001",
"10001111000010011001000010010001",
"00010000000100010101010110001111",
"00001011010100100001000100001111",
"01000010111110001010000000111110",
"00010000000100010000000000100000",
"00111110000100000001000110001001",
"10010000100100011111011110000011",
"00001110000110000000101101010010",
"00101010100100000000110001010001",
"11111100001111101000100000010000",
"11111001101011000011111011110101",
"01000000111110001011000100111110",
"00001000100100001111111111010110",
"00010000000100010000101010010001",
"10001001100010010000100010001001",
"00111101111110001010000100111110",
"01000101010001100000000000000110",
"00110001010011010101000001011000",
"11110000000000000000000000001101",
"10001111001111100101011000111111",
"11111111010100010011111011111000",
"01000110000000000000001100111101",
"01001000001111100100111001001100",
"01101011101100010000110111111111",
"00010111000011010100000000000010",
"00111110101110111011010101010101",
"00000101001111011111100101101110",
"01001110010011000100011000000000"
)
,(
"00001111000011110011000101010000",
"00100100001111100000111100001111",
"11110101100110000011111011110111",
"10010001000010011001000010010001",
"00010001010101100000100110010000",
"01010010000100010000111100010000",
"11111000001000110011111000001011",
"00010001000000000010001001000010",
"00010000000100011000100100010000",
"01010010111101110000011000111110",
"01010001000011100001100000001011",
"00011000000011100001101000001100",
"00111110111100100000001000111110",
"00101111001111101111010101111111",
"00111110100100001001000111111001",
"11010100010000001111100000110010",
"10010001000010001001000011111111",
"10001001000100000001000100001010",
"00111101100010011000100100001000",
"01001100010001100000000000000100",
"10000011001111100100011101001111",
"00001101100100001001000111111110",
"00111111111100000000000000000000",
"10001001000100000001000101010110",
"00111110111110010000010100111110",
"00000000000011011111100011110111",
"01010110010000000000000000000000",
"00111101111110001111100100111110",
"01010011010001100000000000000100",
"10010000100100010100111001001001",
"00010001111111111000011100111110",
"11100000001111101000100100010000",
"00000000000001010011110111111101",
"01001110010010010101001101000110",
"00001101000010001001000001001000",
"01111111111111111111111111111111",
"10010001100010000001000000011100",
"00010001010101100000100110010000",
"00000000000000000000110100010000",
"00111110010101100100000000000000",
"00001111000011111111100011000110",
"10000100001111100000111100001111",
"00111110000100000001000111110110",
"00001011010100111111100010101111",
"00000000000011010000101101010011",
"01010110010000000000000000000000",
"00111110111101100111001000111110",
"00111110100100011111100010101010",
"00010000000011111111100010011011",
"00011000000010110101001010001000",
"00111110000011000101000100001110",
"01000010000111111111011101110001",
"00001000100100001111111111010000",
"00010000000100010000101010010001",
"00111101100010010000100010001001",
"01010011010001100000000000000111",
"01001111010000110100111001001001",
"11111111100011100011111001010011",
"00111101111110000111110100111110",
"01010011010001100000000000000101",
"00111110010101000101001001010001",
"10010000100100011111110111100010",
"11110000000000000000000000001101",
"00010000000100010101011000111111",
"10010001111110000110010100111110",
"11111000010101010011111010010000",
"00010001100010010001000000010001",
"01011111001111101000100100010000",
"11111000010101000011111011110111",
"01000110000000000000010000111101",
"10010001010011100100000101010100",
"00111100001111100000100110010000",
"00001101000010001001000011111000",
"01111111111111111111111111111111",
"00001111100010000001000000011100",
"00010001001011000010001000001111",
"00010001000010101001000110001010",
"00001111111110000010011000111110",
"00001111001101100010001000011010",
"00010000000010100001110000101010",
"00000101001111010010001010001001",
"01000001010101000100011000000000",
"01000100001111100100100001001110",
"01000010001010010000111000000010",
"00001101001000010000000000000001",
"00000010111111111111111111000000",
"01000010001110000001011100000010",
"00101110010001100000000000010000",
"10000100001111100101010100000000",
"00000001000011010011111000000001",
"01000000000000011011110000111110",
"01000010001010010000000000101101",
"01000000110001100000000000011101",
"00100001100001101000111000001000",
"00001001100100001001000101010110",
"01010110000000000011000001000110",
"10011000000000010110011000111110",
"11000010100111111011100010101101",
"10001111100010011111111111110010",
"01000110010101101000100010000101",
"00011000000011110000000000101110",
"00001000000000010101001000111110",
"01000110000000001101101000111110",
"00001110000111100000100001000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000000000000100011110100100010",
"10011001001111100111111001000110",
"11101110101111000011111011111111",
"01000110000000000000001100111101",
"11010100001111100010111000101110",
"00000000101101010011111000000001",
"01000110000000001101110000111110",
"00111110010101010000000000101110",
"01011010001111100000000100011111",
"00001000010000000100011000000001",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111101001000100000010000011001",
"00101110010001100000000000000010",
"00111110111111111101011100111110",
"00000100001111011110111010001010",
"00101110010100110100011000000000",
"00000001101000010011111000101110",
"00111110000000001000001000111110",
"10010000000011100000000010101001",
"01010011100010000001000000101010",
"00001000111100000001100000111110",
"00101110010001100001011110010000",
"00011000100010000001000000000000",
"00111110000000001101111000111110",
"01000000010001100000000100011001",
"00011001000011100001111000001000",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"01000110000000000000001100111101",
"11001000001111100010111001010011",
"11101110010010000011111011111111",
"01000110000000000000010000111101",
"00001101001011100010111001000101",
"00000010111111111111111111000000",
"00101101000000000100000001000110",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"00101010001011010101001100001000",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"00000000000000110011110100000001",
"01000110001011100100010101000110",
"00011000000001100000100001000000",
"01000000010001100001100010010000",
"00010000000000110001011000001000",
"00001000010000000100011010001000",
"00000000000011010011110100000101",
"00101101010101000100010101010011",
"01000011010001010101001001010000",
"01001111010010010101001101001001",
"00001000010000001100011001001110",
"00011001000011100001111000010000",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00011001000101100000111100001111",
"00000000001100000100011000000100",
"01010101000011110010110000010111",
"01000010000111000011100000010111",
"01000000000110010000000000000100",
"00000101000100001111111111101010",
"11000110001111011000100000001000",
"00001000100100000000100001000000",
"00011001000011100001111000010001",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00110000010001100000010000001111",
"00001111001011000001011100000000",
"00011100001110000001011101010101",
"10011001000000000010010001000010",
"00011000000011111001000000011001",
"10001000000100000001100100001110",
"00001001100100001001000101010110",
"00001111000000000000100101000000",
"00001111000001000001011000010000",
"10011000000000110001011000010000",
"11000010100111111011100010101101",
"00001001100010011111111111110001",
"00010001111111111100110101000000",
"10001001000100000000100000000101",
"00001000010000001100011000111101",
"10000100100110011000111010011110",
"10011001100011111010000011001110",
"00010001101000101000010010011001",
"00000000001011010100011000000100",
"00010001000101110010110000010111",
"10010110100011111000111100010110",
"00010000000100010000100010010000",
"00001001100100001001000110001000",
"00010000000000000000011101000000",
"00010000000000111000010010001110",
"10111000101011011001100010001000",
"11111111111100111100001010011111",
"10001000000000110001000010001001",
"10011001100110011000111110011000",
"01000110001111011000100010000101",
"00100110001111100000000001000101",
"00000111010000100010100111111111",
"00101101010001100010000100000000",
"00000000000000110100000000000000",
"00111110000000000010101101000110",
"00000001001111101111111100010101",
"11100100000011010011110100000000",
"00000010000000101111111111111111",
"00110101111011110011100000111110",
"00111110000000000000011001000010",
"00000001010000001111111111110000",
"00000001001111100000100000000000",
"00101101010011010011110100000000",
"00000110010000100000101000111000",
"00000000010101110100011000000000",
"01000110000000000000001101000000",
"00111110000101100000000000110000",
"10010000001111011111111011100101",
"11110101111101000011111010010001",
"10010110001111100000111100001111",
"00111110000011110000111111111000",
"10010000000010101111100000000000",
"11110101110110010011111000001000",
"10010001000100011000101000010001",
"00010000111100111010001000111110",
"10001001000100000001000110001000",
"01000000010001100101011000111101",
"00101010000011110000010100001000",
"01000110000000000000100101000010",
"10110010001111100000000000101101",
"11110010000000000011111011111110",
"00000000000000000000110100001111",
"01000010000111000111111111110000",
"00001111000011110000000000001000",
"01000000111110111000001000111110",
"00001110010101100000000000000010",
"11111111111111111110010000001101",
"00101010100100000000001000000010",
"11110000001111101000100000010000",
"00111110100100001001000111110001",
"10011011001111101111101101101011",
"11110111101011100011111011110101",
"00001010100100010001000100001010",
"11000000000011010001000000010001",
"00000010000000101111111111111111",
"11110010001000100011111000010111",
"00010000111101001000110100111110",
"00001010100100010001000110001000",
"00010101001111100001000000010001",
"11111111011111110011111011110010",
"00000000000001000100001000101011",
"00000000000001000100000010011001",
"11111111010111100011111000001110",
"10001010000100011000101000010001",
"00110110000010011001000110010000",
"11111111111111111100000000001101",
"00010001000101100000001000000010",
"00010000000100010000101010010001",
"01010110000110001000100110001000",
"01000000000010011001000010010001",
"10010000100100010000000000001111",
"00111110111101010100100100111110",
"00110101001111101111111101001101",
"10001001000100000001000111111111",
"10011111101110001010110110011000",
"10001001111111111110101111000010",
"00010000000010010000100100001001",
"11111111111001001000110110001000",
"01000110100000100000001011111111",
"00001110000111100000100001000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"10010001100100000001100100100010",
"00011001000011110000111100001111",
"00010110000010000000010100011001",
"00000000001011011100011010000100",
"00001110100101101010110010010111",
"00000000010000010100011000000100",
"01000010000010100010101000101101",
"00110000010001100000000000000110",
"00000000000000110100000000000000",
"00010111000000000011011101000110",
"00101010000101110001000100011010",
"00110110000100000000111000011111",
"00000000001111110100001000011100",
"00000100000011100001100100001000",
"00101101000000000100000101000110",
"00000110010000100000101000101010",
"00000000001100000100011000000000",
"01000110000000000000001101000000",
"00011000000101110000000000110111",
"00101001000101110001000100001110",
"00001000000000000000010101000010",
"00000000000000100100000011010110",
"00101101010011001101011100001010",
"00000110010000100000101000101010",
"00000000001100000100011000000000",
"01000110000000000000001101000000",
"00001111000101100000000000110111",
"10011001100010000001000000000011",
"10001001111111111011101001000000",
"00000000000010000100001000001010",
"01010110000000000011000101000110",
"00011000111111100010001000111110",
"00001000010000000100011000111101",
"00010110000000010000000001000110",
"00000001000010101010100001000110",
"00001010101010000100011000111101",
"01000110000011100001100100000010",
"00000011000000010000101010101000",
"00111100000000000000001000111101",
"00000110010000100010101000100011",
"00000000001011010100011000000000",
"00111101111111111110011000111110",
"01001111010010000000000000000100",
"11100100000011010100010001001100",
"00000010000000101111111111111111",
"10010000111011001100010000111110",
"00010001000010101001000100001000",
"00101101010011001000100100010000",
"00000000000001110100001000101010",
"00000000001100000100011000001000",
"00010111000000000000010001000000",
"00010110000000000100000101000110",
"00111101111111111011101000111110",
"01001001010100110000000000000100",
"11010001001111100100111001000111",
"00100010000011110000111111111111",
"11111111111101100100001000101100",
"00100011000000000000000100111101",
"00001010101010000100011000001001",
"00001000010000000100011000000010",
"00010110000000010000000001000110",
"00000010001111010001011100001111",
"10010000010100110010001100000000",
"10000000001111100000100110010001",
"11111111110101100011111011111111",
"11111111100101010011111000010001",
"00001010111111111101110100111110",
"00100001000101111000100100010000",
"00001001100100001001000101010110",
"01000110000000000000011101000000",
"01110000001111100000000000100000",
"10111000101011011001100011111111",
"11111111111100111100001010011111",
"00000000000000100011110110001001",
"10010001100100000011111000100011",
"00010001000100000101011000001001",
"00000000011111100011111010001001",
"11111111111100100011111000111101",
"00111101111010101110110100111110",
"00101110010101010000000000000100",
"00111110010101100101001000101110",
"00000011001111011111111111101111",
"01010010001011100101010100000000",
"00001110000010001001000110010000",
"01000010001010010001000000010111",
"00010001001000010000000000000001",
"10011110001111101000100100010000",
"00111110000011100101011011111111",
"00000010001111011111111110000110",
"00111110001011100101010100000000",
"10111011001111101111111111100010",
"00000000000000110011110111101010",
"01010110010100100010111000101110",
"00111101111111111111000000111110",
"01010010001011100000000000000010",
"00000000001001010011111001010110",
"00101110000000000000000100111101",
"00001111100100010000100010010000",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"10001001000100000001000110001000",
"01010110111111110110000000111110",
"11111111010010000011111000001110",
"01000100000000000000001000111101",
"11111111110111000011111000101110",
"00111101111010100111110100111110",
"00101110010001000000000000000100",
"00111110010101100101001000101110",
"00001110010101101111111101000101",
"00111101111111110010110100111110",
"00101110010001000000000000000011",
"10011110001111100100001101010010",
"01000110000011100100010011101001",
"00111101000000011111111111011000",
"01000100010101010000000000000101",
"01000011010100100010111000101110",
"00000010111111111110110001000110",
"00011100000000000001001001000110",
"00010111000000000001001001000110",
"00000001101110110100001000101100",
"00000010111111111110000001000110",
"00000001000000000100011000001110",
"00011000000011100010101000010111",
"00010000000010100101110011000110",
"10001000000100000001011000000010",
"00001010010011000100011000000001",
"01010110000111000010110000000100",
"00000011000010100100110001000110",
"00001110000000010101001101000010",
"00000000000000010000000011000110",
"00101101000000001111111101000110",
"00001000010000100000101000101100",
"01000000010101110000100000000000",
"00111100010000001101100111010010",
"11111110010001100000000000000001",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000001001010010100000000010000",
"00000000111111010100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000010001011001000000",
"00101101000000001111110001000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000100000011",
"00101100001011010000000011111011",
"00000000000011110100001000001010",
"11011000010001100000111000001000",
"11110110000011010000000111111111",
"10111101000001000000000000001110",
"00000000000000001110101001000000",
"00101101000000001111101001000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000011010111",
"00101100001011010000000011111001",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"11000100010000000001000000000001",
"11111000010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000000101100010100000000010000",
"00000000111101110100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000001001111001000000",
"00101101000000001111011001000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000010001011",
"00101100001011010000000011110101",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"01111000010000000001000000000001",
"11110100010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000000011001010100000000010000",
"00000000111100110100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000000101001001000000",
"00101101000000000001101101000110",
"00001001010000100000101000101100",
"01001100010001100000100000000000",
"01000000000100000000001100001010",
"01000110000000000000000000111111",
"00101100001011010000000000011010",
"00000000000011100100001000001010",
"00001010010011010100011000001000",
"01001110010001100101011000000011",
"01000000000100000000001100001010",
"01000110000000000000000000100111",
"00101100001011010000000000011001",
"00000000000011100100001000001010",
"00001010010011010100011000001000",
"01001110010001100101011000000011",
"01000000000100000000001100001010",
"00001110000010000000000000001111",
"00010111000000000001000001000110",
"00000000000001010100001000101010",
"00000011000010100100111001000110",
"01000110000011101000100000010000",
"00101010000101110000000100000000",
"01000110000000000011100001000010",
"00011010000001000000101001001110",
"01000110000110100001101000011010",
"10010000000101100000100101000000",
"10011101100011100000001000011101",
"00010000100111011000111010011101",
"01000010010111000010110100000010",
"00011000000011100000000000011010",
"00010000000000011000100000010000",
"01011100001011010001011000000010",
"00000000000000110100001000011111",
"00001010000011100010000100010111",
"00000011000101100000001000010001",
"00001110000011100000111010001110",
"00001000000010011000100010001001",
"01000100111111100011010101000000",
"11111111110110000100011000001110",
"11010100110001100011110100000001",
"01000110010101111000001011111111",
"10010000000000011111111111100100",
"10010111110011100000100110010001",
"00000000000100001100011010101100"
)
,(
"01010100000000001101011010011100",
"01000010000010100010110000101101",
"10011110000010000000000000000101",
"00000000000000000000111001000000",
"00001010001011000010110101010101",
"00001000000000000000010101000010",
"00000000000000010100000010011000",
"00000000110100101010001000001000",
"00001010001011000010110101010010",
"00001000000000000000011001000010",
"00001110010000001001011110001110",
"00101101010100110000000000000000",
"00000101010000100000101000101100",
"01000000100110100000100000000000",
"10100010000010000000000000000001",
"10000001111111111110010011000110",
"00010110000100000000001001011010",
"00111110000110101000100000010000",
"11101000010001101110101001001000",
"11010100110001100000000111111111",
"11000110001111011000000111111111",
"00010000100000101111111111100100",
"01010110000000000001110001001010",
"01000010000010100010110000101101",
"01010010000010000000000000000101",
"00000000000000000000111101000000",
"00001010001011000010110101001110",
"00001000000000000000010101000010",
"00000000000000100100000001010011",
"01010011000100000101010000001000",
"00101101010101000000000000011100",
"00000101010000100000101000101100",
"01000000010101000000100000000000",
"01010101000000000000000000001111",
"01000010000010100010110000101101",
"01010101000010000000000000000101",
"00001000000000000000001001000000",
"00010000110001100100111101010110",
"00000001110000101001110000000000",
"00000010010110100001100000000000",
"10000010111111111110100011000110",
"10001000000100000001011000010000",
"11101001111001100011111000011010",
"01010011000000000000011000111101",
"01001001010100110101010001000101",
"01010100001111100100111101001111",
"00000100100100000000100100001001",
"10011000000001000001000010011000",
"00010000100110000000010000010000",
"00000100000100001001100000000100",
"10011000001000100010000001001110",
"00010000010001100000010000010000",
"10011000001000100010000000000000",
"01000110000001001000100000010000",
"00100010001000000000000000011000",
"00111101111111110000111100111110",
"01000101010001110000000000000110",
"01001111010010010101001101010100",
"00000110001000010011111001010101",
"00111110000000000001000001000110",
"01001100010001101110011100001000",
"00000000010001100000001000001001",
"00001110000101110000111100000100",
"01001110111001110100010000111110",
"11100111001111110011111000100011",
"11100111001110110011111001010110",
"00111110000000000001101001000110",
"00111110010101111110011011101100",
"01010101001111010000010111111011",
"01000110000001011111011000111110",
"00101100000000100000100101001100",
"01000110000000000011000001000010",
"11010101001111100000000000010000",
"00000100000000000100011011100110",
"11100111000101110011111000001110",
"00010010001111100010001101001110",
"00001110001111100101011111100111",
"00000000000110100100011011100111",
"01000110111001101011111100111110",
"01010101000000101111111111010100",
"00000001111111111101010001000110",
"00000010000010010100110001000110",
"01000110111111111111100101000010",
"01000110000000011111111111010100",
"01000110000000101111111111010100",
"01000110000000100000100101000000",
"00010110000000100000100101001000",
"00001001010011000100011000000100",
"01010110000101110101010100000010",
"00001001010011000100011000100101",
"00001001010010000100011000000001",
"11111111010001100001100000000010",
"01001000010001100001110000000011",
"00001010100100010000000100001001",
"11010100010001101000100000010000",
"00111110010101110000000111111111",
"00000100001111010000010110001011",
"01011001010001010100101100000000",
"10000000001111100101010100111111",
"00101100001011010000111000000101",
"00001000000000000000011101000010",
"01000000111111110111110000111110",
"11111100100011011111111111110100",
"10000010000000101111111111111111",
"10011100110110101001011011010011",
"00110110001011011001111010001110",
"00010000000000000000100101000010",
"01100010001111101001100000000011",
"11111111111100100100000011111111",
"10011001100101111000111100001001",
"00010000100001011000111110011001",
"01001100001111100101011110001000",
"00000000000000110011110100000101",
"00111110010110010100010101001011",
"00001110000111101111111110111111",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000000000001000011110100100010",
"01000100010100100100111101010111",
"11111111110101001100011000001000",
"00001001010010000100011010000010",
"00001001010011000100011000000001",
"11111111110101001100011000000001",
"00000000000001010011110110000001",
"01010011010100100100000101010000",
"11111111110101001100011001000101",
"00001001010011000100011010000010",
"00001001010010000100011000000010",
"11010100110001100101010100000010",
"00001101001111011000000111111111",
"01010011010001010101001000000000",
"01000101010100100100111101010100",
"01010000010011100100100100101101",
"00001110010101100101010001010101",
"11111111110000000011111001010101",
"01010011000000000000101000111101",
"00101101010001010101011001000001",
"01010101010100000100111001001001",
"11111111111010100011111001010100",
"00111101111111101011100100111110",
"01010101010100010000000000000101",
"01010100010110010101001001000101",
"10010000000001001101001000111110",
"11010010001111101101011000001000",
"00111110100100000000111011111110",
"00000011000011111110011001000000",
"10101100100101111100111010001110",
"10001000000000000000111111000010",
"11000010100111111010100110011001",
"01000000000110010000000000000100",
"01000000100110000000000000000001",
"11001100000110000000000000001101",
"00000101110000101010110010010111",
"01000000100011101000101000000000",
"10101101100110000000000000000001",
"11001101110000101001111110111000",
"10001001000100010000100011111111",
"00000100100101010011111001011000",
"01010010000000000000011000111101",
"01001100010010010100011001000101",
"10001000001111100101010101001100",
"11111111101011110011111000000100",
"11111111111111111111000000001101",
"00111110010101110000000100000010",
"00000110001111010000010001111011",
"01000011010000110100000100000000",
"10010000010101000101000001000101",
"00000010000011101001000000001000",
"00000010000011100001110100010110",
"00111000001011010001110100010110",
"10010000000000000100001101000010",
"00011000000011100000001010011101",
"00010001000000000000111001000010",
"00011101000100000001000100010110",
"00111110000000101000100000010000",
"00101010010000000000000000111011",
"00111110000100000000100000000000",
"10001110100111101110001011111011",
"10100000110011101000010010011001",
"10000100100110011001100110001111",
"10010110110100111001011010100010",
"00001001010000101001110011011010",
"00010000000100010000111000000000",
"00111110100100010001000110001000",
"00010000000010000000000001001100",
"00011000000000101000100000010000",
"01000000000101100001101000011010",
"10001001000010011111111110111000",
"01000101000000000000011000111101",
"01000011010001010101000001011000",
"10010000100100010101011001010100",
"00000000001001000100000000001001",
"10010001000000101001110110010000",
"00000011100100001001000100010110",
"10011000001000110100111000010001",
"01000110000100010000001100010000",
"10011000001000110000000000010000",
"01000110000100010000001100010000",
"10011000001000110000000000011000",
"10001001000100010000001100010000",
"10011000100010010001000100010000",
"11000010100111111011100010101101",
"00001010100010011111111111010110",
"00001000100100000011110100001010",
"10011001000100001000001010010000",
"00011101000000001001101001000010",
"00011000000011100000001000001110",
"11111111000011010000111100110110",
"00011100011111111111111111111111",
"00011111001010100001011100010001",
"00000000100000010100001000011100",
"00010110000011110000101010010001",
"00100011010101010001101010010000",
"11000110100001001001000000011001",
"00010001100111000000000010000000",
"10101010000010001001000010001010",
"01001001000000000011000011000010",
"00000010000111010000101101010011",
"00011100000000001111111101000110",
"00101100001011010101001100000000",
"00000000000010000100001000001010",
"00111111010001100000100000001000",
"00000000000011110100000000000000",
"00101100001011010101001000000000",
"00000000000001010100001000001010",
"00000010010000001001111000001000",
"00010000100110000000100000000000",
"00011100000000001000000001000110",
"00011000000000110000111100100010",
"00011101000111010000101101010100",
"00000001010000100100001110011011",
"10010001100100000000001000000000",
"00000011000100000001000100001001",
"10011000001000110100111000010001",
"01000110000100010000001100010000",
"10011000001000110000000000010000",
"01000110000100010000001100010000",
"10011000001000110000000000011000",
"00010001100010100000001100010000",
"00000101010000100001110001010101",
"00010000000110100001000100000000",
"01010111100010010000001100011000",
"10001000000100000000000100010000",
"01100001010000000000100000001110",
"10001001000010010000100011111111",
"01010110000000100000111000111101",
"01000000000010011001000010010001",
"10010000000111010000000000011010",
"11111111000011010001100000000010",
"00011100011111111111111111111111",
"00001010000111110011100000101101",
"00000000000001000100001000001110",
"00111101100010011000100000001010",
"10011000100010000001000000001000",
"11000010100111111011100010101101",
"00001001100010011111111111100000",
"10010000100100010011110101010110",
"00000010000011101001000000001001",
"00000010000011100001110100010110",
"00111000001011010001110100010110",
"10010000000000001000001001000010",
"10101100100101111101011110000010",
"00000000011100001100001000011101",
"00011001000011100001111000001110",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"01011010000101100101001100010110",
"00010001100010000001000000011100",
"00111110000011110000101010010001",
"01010010010000101111111110011111",
"00001110000111100000111100000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11100100001010000011111000100010",
"00000000001011001001101000001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110111001000001010100111110",
"00101010000100011110010001111111",
"01000111000000000010001101000010",
"01000110111000111001001100111110",
"11010110001111100000000000011000",
"01001111001111100001000011100011",
"10010111100100011001000000000110",
"00011000000000100000111100001111",
"10001000000100000001101000011010",
"11100011110110010011111000010110",
"00111110000000000001101001000110",
"10001000000100001110001101110100",
"00001010000010001001000010011000",
"00011010000110000000001000001110",
"01111001010000000001011000011010",
"00010000100010000000100111111111",
"00000000000010100011110110001001",
"01100100011011100111010100100000",
"01101110011010010110011001100101",
"01000110010101010110010001100101",
"10111101000000011111111111010100",
"11111111111111111100110000001101",
"01000110000011100000001000000010",
"00011001000000100000101001111100",
"00010000000010101001000100010110",
"00000010000011100000111010001000",
"10010000000111010001011000011101",
"00010000000011110000111100001000",
"11001110001111100001011100001111",
"00010111000011110001000011111101",
"11111111001011100011111001010110",
"00000000010110000100001000101011",
"11000110100010000001000000001000",
"00111110100000101111111111010100",
"11010100110001101111111111000100",
"00101100000001111000000111111111",
"00001101000000000010011001000010",
"00000010111111111111111111001100",
"01111100010001100000111000000010",
"00010110000110010000001000001010",
"10001000000100000000101010010001",
"00011010010101010000111100001111",
"11111101100101110011111000011010",
"01000110000110100001101001010101",
"00111110000000100000101010000000",
"00011100010000001111111011110100",
"11100011110010010011111000000000",
"00000000001011010011001000001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110111000110100100100111110",
"11001001001111101110001110110011",
"00000000000000010100000011100001",
"00000000010011110011110110001000",
"00101010001010100010101000101010",
"00101010001010100010101000101010",
"01110100011000010110010000100000",
"01110100011100110010000001100001",
"00100000011010110110001101100001",
"01110010011100100110111101100011",
"01100101011101000111000001110101",
"01101000011101000010000001100100",
"01100111011101010110111101110010",
"01101110011010010010000001101000",
"01100001011010010111010001101001",
"01101111011000110010000001101100",
"00100000001011000110010101100100",
"01100011011100100110111101100110",
"01100001001000000111001101100101",
"01110011011001010111001000100000",
"01110100011100100110000101110100",
"00101010001000000010000100100000",
"00101010001010100010101000101010",
"00001101001010100010101000101010",
"00000010111111111111111111001100",
"00001010100001000100011000000010",
"10000000010001100010110000000010",
"00100010001011000000001000001010",
"00001101000000000000111101000010",
"00000010111111111111111111111100",
"00001010011101000100011000000010",
"10000100010001100000111000000001",
"01000110010101100000000100001010",
"01010111000000010000101001011100",
"00000011000010100100111101000110",
"00000000111100000100011001010111",
"01000110000001000001000100111110",
"00100010000000100000101001011100",
"00001010011111000100011000001111",
"01111000010001100000111000000001",
"00101100000010100000000100001010",
"00001101000000000100111001000010",
"00000010111111111111111111001100",
"00010000010100011001000000000010",
"11011111000101000011111000011101",
"00111000111111101101000100111110",
"01000110000100010001111110010000",
"00011001000000100000101001111100",
"01000010000111000000010000010110",
"00001110000100010000000000010010",
"01010010001101010000001010001001",
"00001101000101100001011000011100",
"00000010111111111111111111001100",
"00000000000111010100000000000001",
"10000001000010100111100011000110",
"00000010000010100111010001000110",
"11111111111111111111110000001101",
"01010110100010000000000100000010",
"00001110000010101000010001000110",
"10101100001111100001110100000010",
"11100000000000000011111011011111",
"11011101001111100100011100000001",
"00000000000101000100011011100001",
"01000110111000100010000000111110",
"00111110000000100000101001011100",
"01111000010001100000010010010110",
"01000110001101100000001000001010",
"00111110000101100000000000011010",
"01000110010101101110000111000100",
"00111101000000110000101001001111",
"00000011110011010011111001010111",
"01100001010000100010110010010000",
"00010000000101101001000100000000",
"01000010001110000010110110001000",
"10000010100100000000000001011000",
"00001110000111100000111000011101",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00010110010100110001011000100010",
"00111110000011110001110001011010",
"00001011010000101101111101011011",
"00010000000100011001000100000000",
"10111101001111100101001010001001",
"00000000001010000100000011111100",
"00001111100110001000100000001000",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"11100001000011011110000111101010",
"00011110000001000000000000101110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"11010111001111100010001000000100",
"11100010010000010011111011100001",
"00011000000000100000111000001010",
"01000000000101100001101000011010",
"01010110000010011111111110100011",
"10110101000010101000010001000110",
"01000110000000000001001111000010",
"00001101000000100000101001110100",
"00000010111111111111111111111100",
"00011101000000100000111000000001",
"00111110110111110000001000111110",
"01000111000000011101111101010110",
"01000110111000010011001100111110",
"01110110001111100000000000010100",
"00001110100010000001000011100001",
"00110110000000111110110100111110",
"00010110000000000001101001000110",
"11111111110101000100011001010101",
"11100001000110100011111000000001",
"00100000000000000000101100111101",
"01100101011100100110111001110101",
"01110110011011000110111101110011",
"00111101010011100110010001100101",
"00000011001111010010001001010101",
"01010010010010010100010000000000",
"00000000000000110011110101010010",
"01010100010011100100100101000010",
"01010111000000000000001100111101",
"00111101010100000100111100101111",
"00101111010100100000000000000011",
"11111111110101001100011001001111",
"00001010100111000100011010000010",
"00010110000000100000111100001111",
"00001001000000010000111110010000",
"00001010101001001100011010101100",
"00000011110000101001110010000010",
"00000000000010100011111000000000",
"10000001111111111101010011000110",
"01010010000000000000001100111101",
"01011000010001100101011100101111",
"01000010001101010000001000001010",
"01000110010101100000000000001010",
"00001110000000010000101010100100",
"11011110110101000011111001010111",
"00000000000001110011110100001000",
"01001011010000110100111101001100",
"01000110010011110010111101001001",
"01010110000000101111111111010100",
"00001010010011010100011000001110",
"00001010010111000100011000000011",
"11111111110101000100011000000001",
"00001010010011010100011000000001",
"11111000010000100011011000000100",
"11111111110101000100011011111111",
"00001010010011010100011000000010",
"00000000000110100100011000000100",
"01011100010001100010000100010111",
"01010110000101100000001000001010",
"00001010010011010100011000001110",
"00001010010111000100011000000011",
"11010100010001100000111100000001",
"00111101000010100000000111111111",
"10010000100100010101010101001000",
"00001010010100000100011000001001",
"00100000000100000101010100000010",
"00101100000111000000111100001111",
"00100010000000000000100001000010",
"00000001000010100101000001000110",
"00001001001111011000100100010000",
"10011111101110001010110110011000",
"10001001111111111110001011000010",
"00111110010101010011110101010111",
"11010100110001101111111101010111",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01000111111000000011011100111110",
"10010000111000000111110000111110",
"01000110111000000111100000111110",
"00101001001111100000000000011010",
"11111111011110110011111011100000",
"00000000000100110100001000101011",
"10011011100110111001101110011011",
"00011111001000000001000001010101",
"01010000110001100010001001010101",
"00011100000000100001000000001010",
"10001000100010000000000100010000",
"10000001111111111101010011000110",
"11111111000110010011111001010111",
"00010100001111100101010100111101",
"11111111110101001100011011111111",
"11010100010001100101010110000010"
)
,(
"00001000100100000000000111111111",
"00011010111111111000010100111110",
"00100010000110100001101000011010",
"00011101010000100001111100101001",
"00111110010001111001000000000000",
"00111110000100011101111111100100",
"00100110001111101110000000101001",
"11100000001110010011111011100000",
"00111110000000000001101001000110",
"10001001000100001101111111010100",
"01000000111111110010010000111110",
"00001010100010000000000000000100",
"11010100110001100000111000001010",
"00111110010101111000000111111111",
"00001010001111011111111011010011",
"01001111010011000100001100000000",
"01000110001011010100010101010011",
"00111110010001010100110001001001",
"01010101001000101111111010101110",
"00111101111111111010011000111110",
"11111111101000010011111001010110",
"01000011000000000000101100111101",
"01010100010000010100010101010010",
"01001001010001100010110101000101",
"00111110010101010100010101001100",
"11010100110001101111111010100111",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01001000110111111000011100111110",
"00111110110111111100110000111110",
"00011010010001101101111111011111",
"11011111011110100011111000000000",
"11000110111111101100110000111110",
"01010111100000011111111111010100",
"00111101111111101000001000111110",
"01010000010011110000000000001001",
"01000110001011010100111001000101",
"01010101010001010100110001001001",
"11000110111111100111001000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011111010100100011111001000111",
"11011111100101110011111001010000",
"01000110110111111001010000111110",
"01000101001111100000000000011010",
"11111111111111000000110111011111",
"01010011000000100000001011111111",
"01001110000111000101101000010110",
"00111110000000001111000001000110",
"00111110000010000000000011010010",
"00001000100100001111111010000101",
"11111111111111111111110000001101",
"00010110010100110000001000000010",
"00011101100100000001110001011010",
"00000010100010000001000000000010",
"11010100110001101000100000010000",
"00111110010101111000000111111111",
"00001011001111011111111000100111",
"01001100010001010100010000000000",
"00101101010001010101010001000101",
"01000101010011000100100101000110",
"11111110000101010011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"11110101001111100100011100000001",
"00111010001111100100111011011110",
"11011111001101110011111011011111",
"00111110000000000001101001000110",
"11111100000011011101111011101000",
"00000010000000101111111111111111",
"00011100010110100001011001010011",
"00000000111100000100011001001110",
"00001000000000000111010100111110",
"10010000111111100010100000111110",
"11111111111111000000110100001000",
"01010011000000100000001011111111",
"10010000000111000101101000010110",
"10001000000100000000001000011101",
"11000110100010000001000000000010",
"01010111100000011111111111010100",
"00111101111111011100101000111110",
"01001001010001100000000000001101",
"01010000001011010100010101001100",
"01010100010010010101001101001111",
"00001000010011100100111101001001",
"01000110000000000000100100111101",
"00101101010001010100110001001001",
"01000101010110100100100101010011",
"11111101101010010011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"10001001001111100100011100000001",
"11001110001111100100110011011110",
"11011110111000010011111011011110",
"00111110000000000001101001000110",
"11001110001111101101111001111100",
"11111111110101001100011011111101",
"10000100001111100101011110000001",
"00000000000011000011110111111101",
"01001100010000110100111001001001",
"00101101010001010100010001010101",
"01000101010011000100100101000110",
"11110000010001101001000010010001",
"01000000010001100001110000000000",
"00011101100100000001011000001001",
"10011101000000010001000000000001",
"00001111000100000101011010011101",
"00000001000000010001000010011101",
"00111101100010011000100000010000",
"01001110010010010000000000001000",
"01000100010101010100110001000011",
"00011100010001110100010001000101",
"01000000010001100001101000011010",
"00111101000000100001011000001001",
"11111101010000010011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"00111110100100001001000100000001",
"00001000100100001111111110111110",
"11011110000110100011111001000111",
"11011110010111110011111001010100",
"01011010001111101000101000010001",
"00111110100010100001000111011110",
"00011010010001100000000011010010",
"11011110000001100011111000000000",
"10010000111111010101100000111110",
"00010000000000100001000100001000",
"11111111110101001100011010001001",
"00001000001111100101011110000001",
"00000000000001010011110111111101",
"01000011010011110100110001000010",
"11111100001111100101010101001011",
"11111111110101001100011011111100",
"00001101000010001001000010000010",
"00000010111111111111111111111100",
"01011010000101100101001100000010",
"11110000010001100001000000011100",
"11111111011100000011111000000000",
"00111110010001110000100010010000",
"00010110010001101101110111001100",
"11011110000011110011111000000000",
"00111110000000001111000001000110",
"10001010000100011101111000001001",
"01010101000000001000000100111110",
"00000001111111111101010001000110",
"00111110000000000001101001000110",
"00000010001111101101110110110000",
"00001101000010001001000011111101",
"00000010111111111111111111111100",
"01011010000101100101001100000010",
"00010000000000100001000100011100",
"11111111110101001100011010001001",
"10101000001111100101011110000001",
"00000000000010010011110111111100",
"01000100010000010100010101010010",
"01001100010010010100011000101101",
"10011000001111100101010101000101",
"11111111110101001100011011111100",
"11010100010001100101010110000010",
"10010000100100010000000111111111",
"00011100000000001111000001000110",
"00010110000010010100000001000110",
"00010000000000010001110110010000",
"01010110100111011001110100000001",
"00010000100111010000111100010000",
"10001000000100000000000100000001",
"11011101010111100011111001000111",
"11011101101000110011111001010011",
"11011101100111110011111000010000",
"00000000000110000011111000010001",
"00111110000000000001101001000110",
"00111110100010011101110101001100",
"00001000100100001111110010011101",
"11000110100010000001000000000010",
"01010111100000011111111111010100",
"00111101111111000100111000111110",
"11111100010010010011111001010101",
"11011101011110110011111000001110",
"00111110000011100010001101001110",
"00100011010011101101110101110101",
"11011101011011110011111000001110",
"01101010001111100010001101001110",
"00110000001111100101011111011101",
"00000000000010010011110111111100",
"01000100010000010100010101010010",
"01001110010010010100110000101101",
"11111111110101000011111001000101",
"00111101111111111101000100111110",
"11111100000110010011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"11111001001111100100011100000001",
"00111110001111100100111111011100",
"11011101001110110011111011011101",
"01000110111111111101111000111110",
"11101001001111100000000000011010",
"11111100001110110011111011011100",
"10000001111111111101010011000110",
"11111011111100010011111001010111",
"11101100001111100101010100111101",
"11111111110101001100011011111011",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010011011101110011001100",
"00001110001111101101110100010001",
"11111111101100010011111011011101",
"00111110000000000001101001000110",
"00001110001111101101110010111100",
"11111111110101001100011011111100",
"11000100001111100101011110000001",
"00000000000011110011110111111011",
"01001111010100000100010101010010",
"01001001010101000100100101010011",
"01000110001011010100111001001111",
"01010101010001010100110001001001",
"11000110111110111010111000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011100100011100011111001000111",
"00111110000000000001001001000110",
"11100100001111101101110011010001",
"11111111011100010011111011011100",
"00111110000000000001101001000110",
"11001110001111101101110001111100",
"11111111110101001100011011111011",
"10000100001111100101011110000001",
"00000000000010110011110111111011",
"01001001010100110100010101010010",
"01000110001011010100010101011010",
"01010101010001010100110001001001",
"11000110111110110111001000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"00011011000110110001101100011011",
"00111110110111000100111100111110",
"00011010010001101101110010101011",
"11011100010001100011111000000000",
"10000001111111111101010011000110",
"01010000001111100101011101010110",
"00000000000011000011110111111011",
"00101101010101000100010101010011",
"01000101010011000100100101000110",
"01000101010101000100000101000100",
"11111011001111010011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"00011011000110110001101100000001",
"11011100000110100011111000011011",
"01001001110111000111011000111110",
"01001100110111000101110000111110",
"01000110110111000101100000111110",
"00001001001111100000000000011010",
"11111111110101001100011011011100",
"00111110010101110101011010000001",
"00001010001111011111101100010011",
"01001001010100100101011100000000",
"01000110001011010100010101010100",
"01010101010001010100110001001001",
"11000110111110110000001000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011011111000100011111001000111",
"11011100001001110011111001001010",
"01000110110111000011101000111110",
"11010101001111100000000000011010",
"11111111111111000000110111011011",
"01010011000000100000001011111111",
"01010010000111000101101000010110",
"00111110000000001111000001000110",
"00111110000010001111110101100010",
"00001000100100001111101100010101",
"11111111111111111111110000001101",
"00010110010100110000001000000010",
"00010000000000100001110001011010",
"11111111110101001100011010001000",
"10111100001111100101011110000001",
"00000000000010100011110111111010",
"01010100010010010101001001010111",
"01001001010011000010110101000101",
"00111110010101010100010101001110",
"11010100110001101111101010101011",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01000110110110111000101100111110",
"11001110001111100000000000010011",
"11011011111000010011111011011011",
"00111110000000000001101001000110",
"11111100000011011101101101111100",
"00000010000000101111111111111111",
"00011100010110100001011001010011",
"00000000111100000100011001001110",
"00001000111111010000100100111110",
"10010000111110101011110000111110",
"11111111111111001000110100001000",
"11010011100000100000001011111111",
"00010000100111001101101010010110",
"00000010000100000000001000011101",
"11010100110001101000100100010001",
"00111110010101111000000111111111",
"00001011001111011111101001011111",
"01001100010010010100011000000000",
"01010100010100110010110101000101",
"01010011010101010101010001000001",
"00001100001111010101011000001000",
"01010100010001010100011100000000",
"01001100010010010100011000101101",
"01010100010000010100010001000101",
"00111100001111100101010101000101",
"11111111110101001100011011111010",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010010011101101100011100",
"10010000100100011101101101100001",
"01011010001111100000111000001001",
"00100011010011100000111011011011",
"00111110110110110101010000111110",
"00010000000100011101101101100111",
"01001010001111100000111010001001",
"00100011010011100000111011011011",
"00111110110110110100010000111110",
"00011010010001101101101101010111",
"11011010111100100011111000000000",
"11000110111110100100010000111110",
"01010111100000011111111111010100",
"00111101111110011111101000111110",
"01001100010001100000000000001010",
"00101101010010000101001101010101",
"01000101010011000100100101000110",
"11111001111010010011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"11001001001111100100011100000001",
"11011011000011110011111011011010",
"11011011000010110011111000001110",
"00111110001000110100111000001110",
"00011000001111101101101100000101",
"11110000010001101001000111011011",
"11111100010100000011111000000000",
"00011010010001100000100010010000",
"11011010101010100011111000000000",
"00010001111110011111110000111110",
"00010001000010101001000110001010",
"11000110100010010001000000000010",
"01010111100000011111111111010100",
"00111101111110011010101000111110",
"01000101010100100000000000001011",
"01000101010011010100000101001110",
"01001100010010010100011000101101",
"00000000000100000100011001000101",
"00111101111111111010100100111110",
"00111110000000000001000101000110",
"00001101001111011111111110100010",
"01010011010000100100000100000000",
"01010100010101010100110001001111",
"01001001010001100010110101000101",
"00111110010101010100010101001100",
"11010100110001101111100101111011",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01010010110110100101101100111110",
"00001101110110101010000000111110",
"00000011000000000000000000000000",
"11111111111111111101100000001101",
"10010000100100010000001000000010",
"00000000001001010100000000001001",
"00011110000011100000001000010000",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"00001010000111100010001000000100",
"00010000110110101001001000111110",
"00111110010100100000111000011101",
"01010010000111011101101010001011",
"01010011110110101000011000111110",
"00001000100100000001101000011010",
"10011111101110001010110110010110",
"10001001111111111101010111000010",
"00111110000000000001101001000110",
"11010100110001101101101000010100",
"00111110010101111000000111111111",
"00001100001111011111100100011111",
"01010100010011100100010100000000",
"01010011010001010100100101010010",
"01001100010010010100011000101101",
"11111111110101001100011001000101",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010010111101100111110000",
"00011010010001101101101000110101",
"11011001111001100011111000000000",
"10000001111111111101010011000110",
"01010010000000000000111000111101",
"01000100010001000100000101000101",
"01001001010101000100001101001001",
"01010010010000010100111001001111",
"11111111110101001100011001011001",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010100011101100111000100",
"00000110001111101101101000001001",
"11011010000000110011111011011010",
"00111110000000000001101001000110",
"11010100110001101101100110110100",
"00000100001111011000000111111111",
"01000111010000010101000000000000",
"11111111110101001100011001000101",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00010111010001101101100110011100",
"11011001110111110011111000000000",
"01000110110110011101110000111110",
"10001101001111100000000000011010",
"11111111110101001100011011011001",
"00000000000001010011110110000001",
"01011000001011010101010001000001",
"10010000001111100101010101011001",
"11111111110101001100011011111000",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00011100010001101101100101110000",
"11011001101100110011111000000000",
"00111110000000000001101001000110",
"11010100110001101101100101100100",
"00111110010101111000000111111111",
"00001101001111011111100001101111",
"01000001010010000100001100000000",
"01000011010001010100011101001110",
"01010011010100100100000101001000",
"00111110010101010101010001000101",
"11010100110001101111100001011011",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01000110110110010011101100111110",
"01111110001111100000000000011101",
"00000000000110100100011011011001",
"11000110110110010010111100111110",
"01010111100000011111111111010100",
"00111101111110000011101000111110",
"01000100010000010000000000001010",
"01001110010011110100001101000100",
"01000101010011000100111101010011",
"00001001110001010011111000001111",
"00001111000000000010010001000010",
"00000000000011000100001000110101",
"00010000010001100000001000011101",
"00001111000000100001011000000000",
"00110110110101100100110100111110",
"10010000000000000000110001000010",
"01010110000000100001110100001000",
"10001000000100000000001000010110",
"00001000111111111110000001000000",
"00001001000000000000001001000000",
"00000000000010100011110101010110",
"01000011010000100101010101010011",
"01001111010100110100111001001111",
"00111110000011110100010101001100",
"00100000010000100000100110001011",
"00110101000011100000111100000000",
"00001000000000000000011001000010",
"00000000001001000011111000001111",
"00000000000011000100001000101011",
"00000010000111010000100110010001",
"00010000000000100001011001001110",
"11111111111001010100000010001000",
"00000010010000000000101000001010",
"00111101010101100000100100000000",
"01001110010010010000000000001010",
"01001110010000010101010001010011",
"01000110010011110100010101000011",
"10001011001111100000111100001111",
"00100101010000100010101111111111",
"00110101000011110000100000000000",
"00011101000000000000110001000010",
"00000000000100000100011000000010",
"00111110000011110000001000010110",
"01000010001101101101010111011010",
"00001000100100000000000000001100",
"00010110010100100000001000011101",
"01000000100010000001000000000010",
"01000000000010001111111111100000",
"00001010000010100000000000000010",
"01000011000000000000011000111101",
"01010100010101000101001101000001",
"10010000000010001001000001001111",
"00000000000101010100001000110101",
"00010000000011110000001010011101",
"00011100000100010010010000000010",
"00011100001101100000111100110110",
"00011001000000000000011001000010",
"11101101010000001001110110011101",
"01000010000011100000101011111111",
"00010000000010000000000000000100",
"00111101100010010000001000011101",
"10001000000100000000111010010001",
"11111111110100010011111001011010",
"00000000000000110100001000110101",
"00001000101111010000101000001010",
"00000000001110000010110100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110110110001001110100111110",
"00100001000011011110110111100101",
"00011110000001000000000000111000",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"10000111001111100010001000000100",
"01000110000000100001110111011000",
"00000010000101100000000000010000",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"00010101000011011101100001110010"
)
,(
"00011110000001000000000000111000",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"01011111001111100010001000000100",
"11010110111000100011111011011000",
"00100000000000000000101000111101",
"00100000011101000110111101101110",
"01101110011101010110111101100110",
"00100000000000000000101001100100",
"01100011001000000110011001101111",
"01110011011100110110000101101100",
"01100011000000000000110000100000",
"01110100011100110110111001101111",
"01110100011000110111010101110010",
"00001101001000000111001001101111",
"01000001010001010101001100000000",
"00101101010010000100001101010010",
"01001000010101000100010101001101",
"00001000100100000100010001001111",
"01000010100010100001000110010001",
"00001000100100000000000000011101",
"00001000010100010011111000001110",
"00011101000011110011010100011100",
"00000010000101100101001000000010",
"00011100001101100000111100001111",
"00001010000000000000010101000010",
"11111111111011010100000000001010",
"00001111100010000001000000001001",
"00011111000010000011011000111110",
"00001101000000000101100101000010",
"00000100000000000011100110011011",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"00101110001111101101011111100110",
"00111001011110010000110111101101",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11010111110100000011111000100010",
"11101101000101110011111000010000",
"00000000001110000010000100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00010000110101111011100100111110",
"00010000010001100000001000011101",
"00011110000000100001011000000000",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"10100011001111100010001000000100",
"11010110001001100011111011010111",
"00000111110101010011111000001111",
"00001111000000000011001001000010",
"00011111010000100011010111011010",
"00011101000011110000111100000000",
"00000010000101100100101000000010",
"11111110101000010011111000010000",
"00000000000001100100001000110101",
"00001010000010001001000010001001",
"00011101000010000011110100001010",
"00000010000101100101011000000010",
"11111111110111010100000010011011",
"00011101000010001001000000001000",
"00000010000101100100111000000010",
"11000111010000001000100100010000",
"00111001100110110000110111111111",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11010111010101000011111000100010",
"00001101111011001001110000111110",
"00000100000000000011100000100001",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"00011101000100001101011100111110",
"00000000000100000100011000000010",
"00001110000111100000001000010110",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11010111001010000011111000100010",
"00000000001110010110010000001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00010000110101110001010100111110",
"11101100010110110011111010001000",
"00111101110101011001001100111110",
"01101110001000000000000000010011",
"01100110001000000111010001101111",
"01100100011011100111010101101111",
"01100001011010000010000000101100",
"01100101011011000110010001101110",
"00100000000000000010000000100000",
"01110101001000000110011001101111",
"01100110011001010110010001101110",
"01100100011001010110111001101001",
"01101010011000100110111100100000",
"00100000011101000110001101100101",
"01100001001000000111010001100001",
"01100101011100100110010001100100",
"00000111001000000111001101110011",
"01110100011001010110110100000000",
"00100000011001000110111101101000",
"01011000010001010000000000001011",
"01010100010101010100001101000101",
"01000101010011100010110101000101",
"11111111110101001100011001010111",
"01000100010000100011010110000010",
"00001010100101000100011000000000",
"01000110000111011001000000000010",
"00101011000000100000101010001000",
"00001000000000000001000001000010",
"00111110000000111110100001000110",
"01001101000010000000011001111011",
"01000110000011100000000100001111",
"10010000000000010000101010001000",
"00101101000010001000010000111110",
"00010000010000100000101000111000",
"00001111100010000001000000000000",
"00010110000000111110100001000110",
"00001000000001111100011100111110",
"00001010100010000100011010010000",
"00001010100101000100011000000001",
"10001001000100000001000100000001",
"00000001000101100000001000011101",
"11010100110001100000100000001110",
"00001110001111011000000111111111",
"01000101010110000100010100000000",
"01000101010101000101010101000011",
"01010100010001010100110100101101",
"11000110010001000100111101001000",
"00011010100000101111111111010100",
"00001010100100000100011000011010",
"00101010001011010101001000000010",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"10001100010001100001011010010000",
"01000010001010110000001000001010",
"01000110000010000000000000010000",
"00010000001111100000001111101000",
"00001111010011100000100000000110",
"10001100010001100000111000000001",
"00111110100100000000000100001010",
"00111000001011010000100000011001",
"00000000000100000100001000001010",
"01000110000011111000100000010000",
"00111110000101100000001111101000",
"10010000000010000000011101011100",
"00000001000010101000110001000110",
"00000001000010101001000001000110",
"11010100110001101000100100010001",
"00001001001111011000000111111111",
"01001100010000010101001100000000",
"01000001010000110100111101001100",
"11010100110001100100010101010100",
"10001100110001101000001011111111",
"10000010100111011000001000001010",
"00000010000010101001000001000110",
"01000010001110000010110100001111",
"01010110000111010000000000001001",
"00000001000101100001000000001111",
"10001000111111111111001001000000",
"00001010100100000100011000001001",
"11111111110101001100011000000001",
"00000000000010010011110110000001",
"01001100010011000100000101010110",
"01010100010000010100001101001111",
"11111111110101001100011001000101",
"01000110001101100000111110000010",
"00011100000000100000101010011000",
"00001111000000000000110101000010",
"00010111010101010000001000001110",
"00000000000000110100001000101100",
"00001000000000010000111101010100",
"00000010000010101000110001000110",
"00000001000101100000001000011101",
"10000001111111111101010011000110",
"01010011000000000000011100111101",
"01010100010101100101010001000101",
"11010100110001100101000001001111",
"01000110010101101000001011111111",
"01010111000000010000101001101000",
"00000001000010101001100001000110",
"11111111110101000100011001010101",
"10111010001111100101011000000001",
"10000010100100011001000000000010",
"10001001000100000001000100001001",
"00001001100100001001000101010110",
"00011011100100000000001000001110",
"00101100000101110100111000011010",
"00010000000000000100101101000010",
"00000001000011110010001001010100",
"00010000000110000000100010010000",
"00010000000100010000001000011101",
"00011011000001110100110000111110",
"10010000100100010101011000011011",
"00000000001010000100000000001001",
"00011010000110100001000000001111",
"01010101000011110000001000010110",
"00000000000001010100001000011100",
"00011100000000100000111100110101",
"00000010000011110011010100001010",
"00011100001011000001011101010101",
"11000110000000000000101101000010",
"01010100100000101111111111010100",
"11010100110001100000000100001111",
"10011000000010001000000111111111",
"11000010100111111011100010101101",
"00001001100010011111111111010010",
"10001000000100001000100000010000",
"01000010001011000001011101010100",
"00001000100100000000000100000101",
"00000010000111010001000000011000",
"00000010000101100101011000001110",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"01010010000011100000100010000001",
"00001111001101010000001000010110",
"00101100000101110101010100000010",
"00000000000010110100001000011100",
"10000010111111111101010011000110",
"11000110000000010000111101010100",
"00001000100000011111111111010100",
"00000010000101100100111000001110",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"11000110100100000000100010000001",
"10000010100101100000000000010100",
"11111111111111111000110110001110",
"11000010100111000000000000000000",
"01000110000011100000000001100101",
"00000010000101100000000000100000",
"00000000001010000100011000001111",
"00001111001101010000001000010110",
"00110110000101110101001000000010",
"00000000010010110100001000011100",
"10000010111111111101010011000110",
"11000110000000010000111101010010",
"00010000100000011111111111010100",
"00000000111111111111111100001101",
"00111000000110010001110000000000",
"00000000000100000100011000010000",
"00111000000101110101000000100011",
"00000000001010110100001000100010",
"01010110000011110000001000011101",
"01000000000010011001000010010001",
"00000010000011100000000000011010",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"10011000000111010000100010000001",
"11000010100111111011100010101101",
"00001001100010011111111111100000",
"01000110000000000010111001000000",
"00001110000101100000000000011000",
"10010000100100010101011000000010",
"00000000000110100100000000001001",
"00110101000000100000111000011101",
"00010111010101010000001000001111",
"00001011010000100001110000101100",
"11111111110101001100011000000000",
"00000001000011110101010010000010",
"10000001111111111101010011000110",
"10111000101011011001100000001000",
"11111111111000001100001010011111",
"10001001000100010000100010001001",
"10000010111111111101010011000110",
"11000110000000010000111101010010",
"00011101100000011111111111010100",
"10111000101011011001100000011101",
"11111110100101001100001010011111",
"01000010001011000000100010001001",
"00111010001111101111111001111111",
"01010110000000100000111100000001",
"00001110000010011001000010010001",
"00101100000101110101010100000010",
"00001110000000000000010101000010",
"00001000000001001011001000111110",
"10101101100110000001110100011101",
"11101010110000101001111110111000",
"01000110000010011000100111111111",
"00001000000000101111111111010100",
"00001010100110000100011001010110",
"00000001000011110011111000000001",
"10010001010101100000001000001111",
"00000010000011100000100110010000",
"01000010000111000000111101001110",
"00011100010110010000000000000111",
"00001000010000000000000100001111",
"01000010000111000101000000000000",
"00001111010101010000000000000011",
"10011000000111010001110100000001",
"11000010100111111011100010101101",
"00001001100010011111111111100000",
"10000001111111111101010011000110",
"01010110000000000000001000111101",
"11111111110101001100011000100001",
"00000000111101000011111010000010",
"00000110001010100011111010010000",
"11111111111111111111110000001101",
"00010000010101010000001000000010",
"01010011100010000001000000100000",
"00011010000110100001101000010111",
"00000110001011110011111000010110",
"10010000000010100110000001000110",
"00011101100010000001000000000001",
"00000000010010010011111000000001",
"10000001111111111101010011000110",
"01001101000000000000101000111101",
"00100110010010110101001001000001",
"01000101010001010101011101010011",
"00000100001111100101001001010000",
"00111110000000100000100111110101",
"00001000001111011111111110111011",
"01000101010100100100001100000000",
"01001101010001010101010001000001",
"11111111110101001100011001001101",
"00001010011000000100011010000010",
"00000111010000100011010100000010",
"11111100000011010000111000000000",
"00000001000000101111111111111111",
"01000110000011100001011100001110",
"00000001100100000000101001100000",
"00000001000111011000100000010000",
"10000001111111111101010011000110",
"00001010011000000100011000111101",
"00010000000000100001110110010000",
"01000010001101010000001010001000",
"00001111000011110000000000110101",
"10010001000000010001110100011101",
"00100000000100000101010100001110",
"10001000000100000000111000010110",
"00111110000110100001011101010011",
"00001111000011110000000001010001",
"00011101000011110000111100000001",
"00001111010101100000100000000001",
"00011101000011110101011000000001",
"00111110000011110100110000000001",
"00011101000111010000001000111000",
"00111110000000001111111001000110",
"01000110010101100000000000110101",
"00001001000000010000101001101000",
"01010010000000000000100100111101",
"01000001010001010100110001000101",
"01001101010011010100010101010011",
"00001001100100001001000101010110",
"00001111000000000000101101000000",
"00011101000000010000111100000010",
"00010000000111010000100010010000",
"10111000101011011001100010001000",
"11111111111011111100001010011111",
"01000110001111010000100110001001",
"00001110000000100000101001100000",
"01010110001111010001110100011101",
"01000000000010011001000010010001",
"00001111010101100000000000000101",
"10101101100110000001110100000001",
"11110101110000101001111110111000",
"00111101000010001000100111111111",
"11010110000000000010000011000110",
"10011011100101101000111110001111",
"00101101001000000001000001010101",
"00001111010000100000101001011011",
"10010000100010100001000100000000",
"00010001100010000001000000001000",
"00001001100100001001000110001010",
"00000000000000010100000010001000",
"00011000000100000001000110001010",
"01000010000111110011100000010111",
"00010000010101011111111111011010",
"00100001010111000001011100100000",
"00111101100010010001011000010000",
"00001010001010100010110101010001",
"00001000000000000000001001000010",
"00001010011000001100011000111101",
"10010000100000101001110100010000",
"00001110000110011000001000001000",
"00011010001000010001011100010001",
"01010101000100000001101000011010",
"00010110000101100010000000010001",
"00000010000111010000111010010001",
"01010101000101110001000100001110",
"00101100001001000010000000010000",
"00001000000000000001000001000010",
"00010001000011100000001000001110",
"00100000000100000101010100010111",
"00000010010000100010110000100100",
"00001111010101100000100000000000",
"00010000000000100001110110010000",
"00110110000101110000001010001000",
"01000010000111000011011000001111",
"00001110100100010000000000101100",
"11000000001111101000100000010000",
"00010111000100010000111000000010",
"00100100001000000001000001010101",
"00010000010101010001011000010001",
"00100001001111100000111100100000",
"00010111000100010000100000000000",
"00011111001000000001000001010101",
"00001111000101100001000100011100",
"00010111000110100001101001010100",
"01100110001111100001100000010000",
"00001000000010010000111000000010",
"00000101001111011000100110001000",
"01001101010001000100110000000000",
"10010000100100010100001001010011",
"00010000000010100110000011000110",
"00001000100100001000001010011101",
"01000011010000100000111110000010",
"11111111110101000100011000000000",
"00000010000011100000100000000010",
"00001010001110000010110101010011",
"00000000001000000100011000001111",
"00101100000111000010101000010111",
"00001000000000000001101101000010",
"00000010000111010001110100001110",
"00100000000100010101010100010000",
"00010111000100010000111100010110",
"00011010000110100001101000100001",
"10010001000010101001000100010110",
"00010000000000100101001000111110",
"01000110010101011000100100010001",
"10010001000000011111111111010100",
"10100000000010011001000011010101",
"00010000000101111001011000010000",
"11111111101110010100000010001000",
"00010000000100011000100100001001",
"01011111010000100000111110001001",
"11111111110101000100011000000000",
"00000010000011100000100000000010",
"00001010001110000010110101010011",
"00000000001000000100011000001111",
"01000010000111000010101000010111",
"10010001100100000000000000110011",
"00001111000000100001110100001111",
"00110101000000001000010100111110",
"00010001000000000001001001000010",
"00000000101010100011111000001111",
"00001000010000100011010100001010",
"00011101000111011001000000000000",
"00010000000000010001110100001111",
"01000010001101010000101010001000",
"00001111000100000000000000001010",
"00010111010101000001000101010101",
"11111110011100000011111000100000",
"00000101010000001000100100001000",
"00011101000011100000100000000000",
"01000110010101010000001000011101",
"10010001000000011111111111010100",
"10100000000010011001000011010101",
"00010000000101111001011000010000",
"11111111100111010100000010001000",
"11111111110101000100011000001001",
"11000110001111010000100000000010",
"10001110100000100000101001100000",
"10000010100011111101010100010000",
"00000010000011101001011010100000",
"00010111000100000000111100110110",
"00000111010000100001110000101010",
"00011010000110100101010000000000",
"11111111111011100100000000010110",
"00101100000101110001000000001110",
"01010101000000000001011101000010",
"00100000100100000000001000010001",
"11111111000100100011111000001111",
"01010100000100000101010100001110",
"00111010001111100010000000010111",
"00011000100010000001000011111110",
"00111101100010010000000100010001",
"00010000000010100110000011000110",
"00001000100100001000001010011101",
"00010001010101010001000010000010",
"00010001000011110001011000100000",
"00011010100100000010000100010111",
"00010000000101100001101000011010",
"00101100000000100000111100110110",
"00000000000010000100001000011100",
"00010111000110100001101001010100",
"11111111111011110100000010011001",
"10001000000010100000001000011101",
"10011101100100000011110110001001",
"01100000110001101000001010011101",
"10000010100111010001000000001010",
"00001111100000100000100010010000",
"00010000001000000001000101010101",
"00010001100010100001000100010110",
"00011010000110100001101000010111",
"00001111000010101001000100010110",
"00000001010000010011111000001111",
"10001010000100011000101000010001",
"00010000000010011001000010010001",
"00010111100100010001000110001000",
"00000000000101100100001000110110",
"00010110000110100001101001010100",
"00010111000100010000111110011001",
"00100100001000000001000001010101",
"00010000000011110001011000010001",
"01000000000000001110100000111110",
"10010000000010001111111111100001",
"10001001100010010001000000000001",
"00001110000010001001000000111101",
"00101011111111110111110100111110"
)
,(
"00001000000000000000100001000010",
"00001110111110101100111100111110",
"00101011111111110111000100111110",
"00001000000000000000100101000010",
"11111101111001000011111000001110",
"11111111011001000011111000001110",
"00000000000011000100001000110101",
"00001110111111111000101100111110",
"00000000000001000100001000110101",
"00000001000111010000111100010000",
"00111110001111010000101010001000",
"01000010001010110000000000011011",
"01000110000011110000000000000111",
"00000001000011110000000000010000",
"00000000000011010011110100001000",
"01010100010100110100010101000010",
"01000101010001010101001001000110",
"01000011010011110100110001000010",
"01010000010000100011010101001011",
"11111111110101001100011000000000",
"01011010000101100100101110000010",
"01101000010001100000111000011100",
"01000110000101100000001000001010",
"00111110000000010000101001101000",
"11011010001111101111110101100010",
"00010011010000100011010111111110",
"00111110000011110000111100000000",
"01000010001101011111111110001011",
"00011101000111010000000000001001",
"01010101000000010001110100001111",
"00001010000011100000000100001111",
"10001000000100000000101010010001",
"00011100001101100000111100110110",
"00001110000000000001001001000010",
"00001111010101010000001000011101",
"00010111000110100001101001010100",
"00100000000101110101010000000010",
"00010110001111100001011101010100",
"11111111110101001100011011111101",
"00001000001111010010101110000001",
"01001100010011000100000100000000",
"01010100010000010100001101001111",
"01100000001111100101010101000101",
"00001010011000000100011011101110",
"11001111100100000001011100000010",
"00011011000110111010110010011100",
"10011100101110001001000000011011",
"01100100010001100101010100011001",
"00010111010100110000001000001010",
"00010000001010100001011100100000",
"00111110010101110001110010001000",
"00000110001111011110111000111111",
"01001100010000010100110100000000",
"10010000010000110100111101001100",
"10010000100000101001000000001000",
"00001111000011111000001010011101",
"00101100000100010000000100011101",
"00001111000000000000001101000010",
"00010000000010000000000100001111",
"01010110000000010001110100001111",
"01000010000100000000000100001111",
"00010000000011100000000000000011",
"00001000100100001000100100000001",
"00111101100000011001110110011101",
"01000001010010000000000000001011",
"01000101010011000100010001001110",
"01001001010011000100000101010110",
"10010001100000101001000101000100",
"01000010000100001000001010011101",
"00010000000100010000000000000110",
"00000000000000110100000000000001",
"00010001000000010000111100010001",
"00010000000000000000011101000010",
"01000000000000010001110100010001",
"00001111000100000000000000000100",
"00001001100010010000000100011101",
"11111111110101001100011000111101",
"01110000001111100000111010000010",
"00000010000111010000111111111111",
"01000010000011100001110000110110",
"00001000100100000000000001101010",
"11000110000000010000111101010110",
"10011101000100000000101001100000",
"10000010000010001001000010000010",
"10010000000111010000111011010110",
"10000001000101110100111000000010",
"00100000000100010101010100010000",
"00010001000000100000111100010110",
"00011010001000010001011110010001",
"00001111000101100001101000011010",
"00010000010101010001011100010001",
"00010110000100010010010000100000",
"00101101010100110000001000001110",
"01000110000011110000101000111000",
"00101010000101110000000000100000",
"00001111001011000000101000011100",
"00010000000000100001110100011101",
"01000010000111000010110000010111",
"00111110000011110000000000011001",
"00010001000011111111111101111111",
"00100000000100000101010100010111",
"00010110000100010001110000011111",
"00010000000010100000101010010001",
"10011000000101110100111010001000",
"00001000111111111100010001000000",
"00101110001111101000100000010000",
"10001000000100001000100111111111",
"11111111110101001100011000001010",
"00111110000011110011110110000001",
"10011011010000101111111011110011",
"11111111110101001100011000000000",
"01011010000101100101001110000010",
"00000010000111010000111100011100",
"00010111000110100001101001010100",
"00100000000011110101010100000010",
"00001111000010100001011101001110",
"00000100010000100011100000101101",
"00010000000010101001000100000000",
"00000101001111100000100010001000",
"00101101000111000101101000000001",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"10010000000110110001101100001000",
"00000010000111010000111100001000",
"11111111111111111111110000001101",
"01010011100100000000001000000010",
"00010001000111000101101000010110",
"00010110010100110001101000011010",
"00000000000000010001010000111110",
"00111110000100010000000000000000",
"10000010100100011111101110000010",
"00000001000011110101010100001111",
"00001000111111110001111000111110",
"10101011001111100001011001001110",
"00001111000011110000111111111011",
"00110101111111011101101000111110",
"00011101000000000000100101000010",
"00000001000111010000111100011101",
"00001110000000010000111100010000",
"00001010100100011000100000001010",
"00001111001101101000100000010000",
"00001100010000100001110000110110",
"00010110010100110001000000000000",
"00011101000011110001110001011010",
"01000111001111100001000100000010",
"11111111111111001000110111111011",
"10001000100000010000001011111111",
"11111111110101001100011000101100",
"00000000000001000100000010000001",
"11111101110100110011111000001010",
"01000110000000000000010000111101",
"11000110010001010100010101010010",
"00001110100000101111111111010100",
"01000010111111100100001000111110",
"00000010000111010000000000010100",
"00010111000110100001101001010100",
"00001010100100010101010100000010",
"01010100001000001000100000010000",
"01000000000101110001101000011010",
"00010111000011100000000000000010",
"10000001111111111101010011000110",
"01010010000000000000011000111101",
"01011010010010010101001101000101",
"11111111110101001100011001000101",
"00010100001111100000111010000010",
"00000000000001010100001011111110",
"00001111000110000000001000001110",
"11010100110001100000100000000001",
"00001110001111011000000111111111",
"01001100010011000100000100000000",
"01010100010000010100001101001111",
"01010011001011010100010001000101",
"11000110010001010101101001001001",
"00001110100000101111111111010100",
"01000010111111011110111000111110",
"00000010000011100000000000010000",
"01010110100100000001011101010101",
"10101100000000010000111100100101",
"00111110000000000000001111000010",
"11000110000010001111111001100011",
"00111101100000011111111111010100",
"01001110010010010000000000001100",
"01000110010001010101001001000011",
"01001110010001010101001001000101",
"11011000000011010100010101000011",
"00000010000000101111111111111111",
"11111111111111111111110000001101",
"00111101000101110000001000000010",
"01000101010001000000000000001100",
"01000110010001010101001001000011",
"01001110010001010101001001000101",
"11111100000011010100010101000011",
"00000010000000101111111111111111",
"00011100010110100001011001010011",
"11111111111111111111110000001101",
"00000110001111010000000100000010",
"01010101010011100101010100000000",
"00001101010001000100010101010011",
"00000010111111111111111111111100",
"11111100000011010001011000000010",
"00000001000000101111111111111111",
"01000001000000000000010100111101",
"01001110010001110100100101001100",
"11001100110010100011111001000111",
"00111110000000000001010101000110",
"10101001001111101100110100001101",
"11101111100001000011111011111111",
"00001010011001000100011001010101",
"00011010001000000001100100000010",
"00001101111011110111100100111110",
"00000100000000000000000000000000",
"11111111111111111100110000001101",
"00111110000101110000001000000010",
"00011010010001101110111101101010",
"11001100100111100011111000000000",
"01000001000000000000010100111101",
"01010100010011110100110001001100",
"00011100010100110011110101010000",
"01010100000000000001000000111101",
"01000111010001110100100101010010",
"01010011001011010101001001000101",
"01001100010000110101001101011001",
"01010010010010110100001101001111",
"01010100000000000001000100111101",
"01000111010001110100100101010010",
"01010000001011010101001001000101",
"01000011010100110100010101010010",
"01010010010001010100110001000001",
"00000000000011010011110101001111",
"01000111010010010101001001010100",
"00101101010100100100010101000111",
"01010101010100000100111001001001",
"01010011000111000101001101010100",
"01000010000010100010110000101101",
"01000111000010000000000000000101",
"01001100000000000000001001000000",
"00111110000011110000111100010110",
"00001111010101011100101100011010",
"11010000010001100010000000011001",
"01000110001000100000001011111111",
"00001001000000011111111111010000",
"01001100000000000000110000111101",
"00101101010010110100001101001111",
"01001110010101010100111101000011",
"00011010010100100100010101010100",
"00001111001000100001101000011010",
"11000000010001100001101000011010",
"00001000000000010001011011111111",
"01010011000000000001001100111101",
"01000011001011010101010001000101",
"01010100010011100101010101001111",
"01010011001011010101001001000101",
"01001001010101100101001001000101",
"00011010000110100100010101000011",
"00010110111111111100000001000110",
"00000000000010100011110100000010",
"01000011010101000100010101010011",
"01010100010011100101010101001111",
"01000110010000110101001001000101",
"11000110000000101111111111010100",
"10010000000100000000101001101100",
"10001000000100000000001000011101",
"10010001010101010101011000000010",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00000001100100001000100000010000",
"00000001000111011000100000010000",
"11111111110110000100011000001110",
"00001010010101000100011000000001",
"10011000010001100011010100000010",
"00011100001011000000001000001010",
"01000110000000000010000101000010",
"01000110000000100000101001100100",
"01011011001011010000000000100000",
"00000000000001000100001000001010",
"00001010001000000000111101010101",
"01101000010001100010001101010100",
"01011011000101110000001000001010",
"00001110000000000000010101000010",
"11001001101110000011111001010111",
"10100100010001100101010100001000",
"10011100010001100000000100001010",
"01000010001011000000001000001010",
"11000001001111100000000000000011",
"11111111110101000100011011101010",
"00001011001111010100010000000001",
"01000001010001010101001000000000",
"01010101010011110100001101000100",
"01010010010001010101010001001110",
"01010011010101100000000000000110",
"01001011010000110100000101010100",
"01001100010101100000000000000111",
"01010100010001110100111001000101",
"01010011000000000000010101001000",
"01010000010001010100010101010111",
"01011001010100110000000000001000",
"01001111010011000100001101010011",
"00000000000010010100101101000011",
"01010010010101010100111101010011",
"01001001001011010100010101000011",
"00100011000000000000010001000100",
"00000011011000100110100101110100",
"01101110011010010011111000000000",
"01101001011101000000000000000011",
"01001000000000000000001101100010",
"00000000000000110100010001001100",
"00001001010001000100000101010000",
"01010110010000010100101000000000",
"01001101010010010101010001000001",
"00000000000000000101001001000101",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000"
)
                           );
  type dvec is array (0 to 9 - 1) of DataVec;
  signal bdata: dvec;
  signal old: std_ulogic_vector(ROMrange'high downto 11);
  
begin
  
  fetch: process(Clock) is
  begin
    if rising_edge(Clock) then
         old <= Address(old'range);
	   for i in bdata'range loop
	     bData(i) <= ROM(i)(to_integer(std_ulogic_vector(Address(11 - 1 downto 2))) MOD blocks'length);
		end loop;
	 end if;
  end process fetch;

  Data <= 
          bdata(0 ) when unsigned(old) = 0 else
          bdata(1 ) when unsigned(old) = 1 else
          bdata(2 ) when unsigned(old) = 2 else
          bdata(3 ) when unsigned(old) = 3 else
          bdata(4 ) when unsigned(old) = 4 else
          bdata(5 ) when unsigned(old) = 5 else
          bdata(6 ) when unsigned(old) = 6 else
          bdata(7 ) when unsigned(old) = 7 else
          bdata(8 ) when unsigned(old) = 8 else
          (others => '0');
			 
end RTL;
