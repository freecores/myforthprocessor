----------------------------------------------------------------------------------
-- Company: RIIC
-- Engineer: Gerhard Hohner Mat.nr.: 7555111
-- 
-- Create Date:    01/07/2004 
-- Design Name:    Diplomarbeit
-- Module Name:    ROMcode - Rtl 
-- Project Name:   32 bit FORTH processor
-- Target Devices: Spartan 3
-- Tool versions:  ISE 8.2
-- Description: implements a ROM containing the BIOS
-- Dependencies: global.vhd
-- 
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------


library IEEE, work;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use work.global.all;

entity ROMcode is
  port (Clock: in std_ulogic;									-- system clock
        Address: in std_ulogic_vector(ROMrange);		-- address bus
		  Data: out DataVec);									-- outgoing data
end ROMcode;

architecture RTL of ROMcode is
  type blocks is array (0 to 2048 / 4 - 1) of DataVec;
  type myarray is array (natural range <>) of blocks;
  constant ROM: myarray := (
(
"01000110010011100101011001010100",
"10101010001111100010010110000000",
"00000000000110110100011000100110",
"00000001111111111111000001000110",
"00111001000000000001011101000110",
"00000000000110000100011000000001",
"00001110010101100000000100110100",
"10010000000010100110110001000110",
"00011101100010000001000000000001",
"11111101001111100101001100000001",
"01000110000000100101101001000001",
"11110110001111100000001111101000",
"01000010011000010011111000010010",
"00000010111111111101010001000110",
"00100110110111000011111000001000",
"00001101001001100111010000111110",
"00000011000000000000000000000000",
"11111111111111111101100000001101",
"01000110010101100000000100000010",
"01010110000000010000101001000000",
"00000001000010100100010001000110",
"01100000010001100000111001010110",
"00010000000000011001000000001010",
"01010110000000010001110110001000",
"00000001000010101000000001000110",
"00001010100001000100011001010110",
"10011000010001100101011000000001",
"01000110010101100000000100001010",
"01010110000000010000101010010000",
"00000001000010101001010001000110",
"00001010100010000100011001010110",
"10001100010001100101011000000001",
"01000110010101100000000100001010",
"01000110000000010000101001101000",
"00001101010100100000101010101100",
"00000100000000000000110100111110",
"00000000000011000101100100111110",
"01010010010101100000000000000000",
"00000000000011010011100000001101",
"00001100010011000011111000000100",
"01001100000000000000000000000000",
"00001101001100100000110101010010",
"00111111001111100000010000000000",
"00000000000000000000000000001100",
"00000000000000000000000000001101",
"00101001000011010101001000000011",
"00111110000001000000000000001101",
"00000000000000000000110000101110",
"00000000000000000000110100000000",
"00001101010100100000001100000000",
"00000100000000000000110100011110",
"00000000000011000001110100111110",
"00010000010001100000000000000000",
"00010011000011010101001000000000",
"00111110000001000000000000001101",
"00000000000000000000110000001110",
"00001010011011000100011000000000",
"00001101000001010000110101010010",
"11111111001111100000010000000000",
"00000000000000000000000000001011",
"00000000000011001110110000001101",
"01110101000011010101001100000100",
"00111110000001000000000000001101",
"11000001000011010000101111101110",
"01010011000001000000000000001101",
"00000000000011100001001000001101",
"00001011111000000011111000000100",
"00000000000011011100110100001101",
"01110110000011010101001100000100",
"00111110000001000000000000001110",
"00011000000011010000101111010010",
"01010011000001000000000000001110",
"00000000000011101100011100001101",
"00001011110001000011111000000100",
"00000000000011101101000000001101",
"11011100000011010101001100000100",
"00111110000001000000000000001110",
"11010110000011010000101110110110",
"01010011000001000000000000001110",
"00000000000011101110101100001101",
"00001011101010000011111000000100",
"00000000000011101110011100001101",
"00011111000011010101001100000100",
"00111110000001000000000000001111",
"11110110000011010000101110011010",
"01010011000001000000000000001110",
"00000000000011110010100100001101",
"00001011100011000011111000000100",
"00000000000011110010010100001101",
"10100010000011010101001100000100",
"00111110000001000000000000001111",
"11110000000011010000101101111110",
"01010011000001000000000000001111",
"00000000000100000011110000001101",
"00001011011100000011111000000100",
"00000000000100000111000000001101",
"10011100000011010101001100000100",
"00111110000001000000000000010000",
"10000110000011010000101101100010",
"01010011000001000000000000010000",
"00000000000100001100101000001101",
"00001011010101000011111000000100",
"00000000000100001010001000001101",
"11010101000011010101001100000100",
"00111110000001000000000000010000",
"11010000000011010000101101000110",
"01010011000001000000000000010000",
"00000000000100001111100000001101",
"00001011001110000011111000000100",
"00000000000100001101110100001101",
"00010011000011010101001100000100",
"00111110000001000000000000010001",
"11111111000011010000101100101010",
"01010011000001000000000000010000",
"00000000000100010011010000001101",
"00001011000111000011111000000100",
"00000000000100010001011100001101",
"01011101000011010101001100000100",
"00111110000001000000000000010010",
"01100110000011010000101100001110",
"01010011000001000000000000010010",
"00000000000100100111101100001101",
"00001011000000000011111000000100",
"00000000000100100111011000001101",
"10101001000011010101001100000100",
"00111110000001000000000000010010",
"10000011000011010000101011110010",
"01010011000001000000000000010010",
"00000000000100101100011100001101",
"00001010111001000011111000000100",
"00000000000100101011000100001101",
"11110001000011010101001100000100",
"00111110000001000000000000010010",
"11001111000011010000101011010110",
"01010011000001000000000000010010",
"00000000000100110000111100001101",
"00001010110010000011111000000100",
"00000000000100110001001100001101",
"00100100000011010101001100000100",
"00111110000001000000000000010011",
"00011000000011010000101010111010",
"01010011000001000000000000010011",
"00000000000100110010110000001101",
"00001010101011000011111000000100",
"00000000000100110010011100001101",
"00110111000011010101001100000100",
"00111110000001000000000000010011",
"00110010000011010000101010011110",
"01010011000001000000000000010011",
"00000000000100110100010100001101",
"00001010100100000011111000000100",
"00000000000100110011101000001101",
"01001111000011010101001100000100",
"00111110000001000000000000010011",
"01001010000011010000101010000010",
"01010011000001000000000000010011",
"00000000000101000010010000001101",
"00001010011101000011111000000100",
"00000000000100110101011000001101",
"00111000000011010101001100000100",
"00111110000001000000000000010100",
"00101000000011010000101001100110",
"01010011000001000000000000010100",
"00000000000101001001010000001101",
"00001010010110000011111000000100",
"00000000000101000100000100001101",
"11100100000011010101001100000100",
"00111110000001000000000000010100",
"10011101000011010000101001001010",
"01010011000001000000000000010100",
"00000000000101010011001000001101",
"00001010001111000011111000000100",
"00000000000101001110110000001101",
"01110110000011010101001100000100",
"00111110000001000000000000010101",
"00111010000011010000101000101110",
"01010011000001000000000000010101",
"00000000000101011011101100001101",
"00001010001000000011111000000100",
"00000000000101010111111000001101",
"11110111000011010101001100000100",
"00111110000001000000000000010101",
"10111111000011010000101000010010",
"01010011000001000000000000010101",
"00000000000101100000011000001101",
"00001010000001000011111000000100",
"00000000000101011111101100001101",
"01010000000011010101001100000100",
"00111110000001000000000000010110",
"00001100000011010000100111110110",
"01010011000001000000000000010110",
"00000000000101101010100100001101",
"00001001111010000011111000000100",
"00000000000101101010111000001101",
"01100101000011010101001100000100",
"00111110000001000000000000010111",
"01101101000011010000100111011010",
"01010011000001000000000000010111",
"00000000000110001000010100001101",
"00001001110011000011111000000100",
"00000000000110001011101000001101",
"10101110000011010101001100000100",
"00111110000001000000000000011001",
"10100111000011010000100110111110",
"01010011000001000000000000011001",
"00000000000110011011100100001101",
"00001001101100000011111000000100",
"00000000000110011011001000001101",
"00100100000011010101001100000100",
"00111110000001000000000000011010",
"10111101000011010000100110100010",
"01010011000001000000000000011001",
"00000000000110101010110100001101",
"00001001100101000011111000000100",
"00000000000110100010100000001101",
"11111011000011010101001100000100",
"00111110000001000000000000011010",
"10111001000011010000100110000110",
"01010011000001000000000000011010",
"00000000000110110010100000001101",
"00001001011110000011111000000100",
"00000000000110110000000000001101",
"01010000000011010101001100000100",
"00111110000001000000000000011011",
"00110000000011010000100101101010",
"01010011000001000000000000011011",
"00000000000110110111011000001101",
"00001001010111000011111000000100",
"00000000000110110101011100001101",
"10100101000011010101001100000100",
"00111110000001000000000000011011",
"01111100000011010000100101001110",
"01010011000001000000000000011011",
"00000000000110111011101100001101",
"00001001010000000011111000000100",
"00000000000110111010101100001101",
"11010111000011010101001100000100",
"00111110000001000000000000011011",
"11000011000011010000100100110010",
"01010011000001000000000000011011",
"00000000000110111111011000001101",
"00001001001001000011111000000100",
"00000000000110111101110000001101",
"00001110000011010101001100000100",
"00111110000001000000000000011100",
"11111101000011010000100100010110",
"01010011000001000000000000011011",
"00000000000111000011001100001101",
"00001001000010000011111000000100",
"00000000000111000001011000001101",
"01010100000011010101001100000100",
"00111110000001000000000000011100",
"00111010000011010000100011111010",
"01010011000001000000000000011100",
"00000000000111001010010100001101",
"00001000111011000011111000000100",
"00000000000111000101101100001101",
"11010101000011010101001100000100",
"00111110000001000000000000011100",
"10101101000011010000100011011110",
"01010011000001000000000000011100",
"00000000000111010000001100001101",
"00001000110100000011111000000100",
"00000000000111001101110000001101",
"01010110000011010101001100000100",
"00111110000001000000000000011101",
"00001011000011010000100011000010",
"01010011000001000000000000011101",
"00000000000111010111110000001101",
"00001000101101000011111000000100",
"00000000000111010101111000001101",
"11000101000011010101001100000100",
"00111110000001000000000000011101",
"10000010000011010000100010100110",
"01010011000001000000000000011101",
"00000000000111011101100100001101",
"00001000100110000011111000000100",
"00000000000111011100110000001101",
"10010000000011010101001100000100",
"00111110000001000000000000011110",
"11011111000011010000100010001010",
"01010011000001000000000000011101",
"00000000000111101010010100001101",
"00001000011111000011111000000100",
"00000000000111101001100000001101",
"10111011000011010101001100000100",
"00111110000001000000000000011110",
"10101010000011010000100001101110",
"01010011000001000000000000011110",
"00000000000111110000110000001101",
"00001000011000000011111000000100",
"00000000000111101100001000001101",
"00110000000011010101001100000100",
"00111110000001000000000000011111",
"00010010000011010000100001010010",
"01010011000001000000000000011111",
"00000000000111110100001000001101",
"00001000010001000011111000000100",
"00000000000111110011011000001101",
"10011100000011010101001100000100",
"00111110000001000000000000011111",
"01001001000011010000100000110110",
"01010011000001000000000000011111",
"00000000000111111010110000001101",
"00001000001010000011111000000100",
"00000000000111111010010100001101",
"11010101000011010101001100000100",
"00111110000001000000000000011111",
"10110011000011010000100000011010",
"01010011000001000000000000011111",
"00000000001000000000001100001101",
"00001000000011000011111000000100",
"00000000000111111101101100001101",
"01101010000011010101001100000100",
"00111110000001000000000000100000",
"00001010000011010000011111111110",
"01010011000001000000000000100000",
"00000000001000000111010100001101",
"00000111111100000011111000000100",
"00000000001000000110111000001101",
"10011100000011010101001100000100",
"00111110000001000000000000100000",
"01111010000011010000011111100010",
"01010011000001000000000000100000",
"00000000001000001010011100001101",
"00000111110101000011111000000100",
"00000000001000001010000000001101",
"11011101000011010101001100000100",
"00111110000001000000000000100000",
"10101101000011010000011111000110",
"01010011000001000000000000100000",
"00000000001000001110100100001101",
"00000111101110000011111000000100",
"00000000001000001110001000001101",
"00001110000011010101001100000100",
"00111110000001000000000000100001",
"11101111000011010000011110101010",
"01010011000001000000000000100000",
"00000000001000010010011000001101",
"00000111100111000011111000000100",
"00000000001000111000111000001101",
"10100110000011010101001100000100",
"00111110000001000000000000100011",
"10011010000011010000011110001110",
"01010011000001000000000000100011",
"00000000001000111011010100001101",
"00000111100000000011111000000100",
"00000000001000111010101000001101",
"11100001000011010101001100000100",
"00111110000001000000000000100011",
"10111011000011010000011101110010",
"01010011000001000000000000100011",
"00000000001000111111001000001101",
"00000111011001000011111000000100",
"00000000001000111110011100001101",
"00000100000011010101001100000100",
"00111110000001000000000000100100",
"11110101000011010000011101010110",
"01010011000001000000000000100011",
"00000000001001000011001100001101",
"00000111010010000011111000000100",
"00000000001001000011011100001101",
"01001001000011010101001100000100",
"00111110000001000000000000100100",
"01000010000011010000011100111010",
"01010011000001000000000000100100",
"00000000001001000101010000001101",
"00000111001011000011111000000100",
"00000000001001000100111100001101",
"01110000000011010101001100000100",
"00111110000001000000000000100100",
"01011001000011010000011100011110",
"01010011000001000000000000100100",
"00000000001001000111101100001101",
"00000111000100000011111000000100",
"00000000001001000111010000001101",
"10000101000011010101001100000100",
"00111110000001000000000000100100",
"10000000000011010000011100000010",
"01010011000001000000000000100100",
"00000000001001001000111000001101",
"00000110111101000011111000000100",
"00000000001001001000100100001101",
"10101110000011010101001100000100",
"00111110000001000000000000100100",
"10010001000011010000011011100110",
"01010011000001000000000000100100",
"00000000001001001011100100001101",
"00000110110110000011111000000100",
"00000000001001001011001000001101",
"11001001000011010101001100000100",
"00111110000001000000000000100100",
"10111111000011010000011011001010",
"01010011000001000000000000100100",
"00000000001001001101100100001101",
"00000110101111000011111000000100",
"00000000001001101011001100001101",
"01110010000011010101001100000100",
"00111110000001000000000000100111",
"00011000000011010000011010101110",
"01010011000001000000000000100111",
"00000000001001111010010100001101",
"00000110101000000011111000000100",
"00000000001001111010110100001101",
"01001000000011010101001100000100",
"00111110000001000000000000101000",
"11011000000011010000011010010010",
"01010011000001000000000000100111",
"00000000001010001000011100001101",
"00000110100001000011111000000100",
"00000000001010000100111000001101",
"10011011000011010101001100000100",
"00111110000001000000000000101000",
"10001100000011010000011001110110",
"01010011000001000000000000101000",
"00000000001010001011001100001101",
"00000110011010000011111000000100",
"00000000001010001010000100001101",
"11001100000011010101001100000100",
"00111110000001000000000000101000",
"10111010000011010000011001011010",
"01010011000001000000000000101000",
"00000000001010001110001000001101",
"00000110010011000011111000000100",
"00000000001010001101101100001101",
"11110101000011010101001100000100",
"00111110000001000000000000101000",
"11101110000011010000011000111110",
"01010011000001000000000000101000",
"00000000001010010011111000001101",
"00000110001100000011111000000100",
"00000000001010001111110000001101",
"01011000000011010101001100000100",
"00111110000001000000000000101001",
"01000110000011010000011000100010",
"01010011000001000000000000101001",
"00000000001010011011011000001101",
"00000110000101000011111000000100",
"00000000001011011011000000001101",
"10110101000011010101001100000100",
"00111110000001000000000000101101",
"10110010000011010000011000000110",
"01010011000001000000000000101101",
"00000000001011011011110000001101",
"00000101111110000011111000000100",
"00000000001011011011101000001101",
"11000011000011010101001100000100",
"00111110000001000000000000101101",
"11000001000011010000010111101010",
"01010011000001000000000000101101",
"00000000001011011100101000001101",
"00000101110111000011111000000100",
"00000000001011011100100000001101",
"11101111000011010101001100000100",
"00111110000001000000000000101101",
"11001111000011010000010111001110",
"01010011000001000000000000101101",
"00000000001011100000100000001101",
"00000101110000000011111000000100",
"00000000001011100111010000001101",
"11111101000011010101001100000100",
"00111110000001000000000000101110",
"00001001000011010000010110110010",
"01010011000001000000000000101111",
"00000000001011110001011100001101",
"00000101101001000011111000000100",
"00000000001011110001001000001101",
"01001110000011010101001100000100",
"00111110000001000000000000101111",
"00100100000011010000010110010110",
"01010011000001000000000000101111",
"00000000001011111010100100001101",
"00000101100010000011111000000100",
"00000000001011110101100100001101",
"00000110000011010101001100000100",
"00111110000001000000000000110000",
"10110110000011010000010101111010",
"01010011000001000000000000101111",
"00000000001100000001011100001101",
"00000101011011000011111000000100",
"00000000001100000001010100001101",
"01001100000011010101001100000100",
"00111110000001000000000000110000",
"00100010000011010000010101011110",
"01010011000001000000000000110000",
"00000000001100000111011000001101",
"00000101010100000011111000000100",
"00000000001100001000000000001101",
"11001000000011010101001100000100",
"00111110000001000000000000110000",
"10001010000011010000010101000010",
"01010011000001000000000000110000",
"00000000001100010010100000001101",
"00000101001101000011111000000100",
"00000000001100010011001100001101",
"10100000000011010101001100000100",
"00111110000001000000000000110001",
"10110010000011010000010100100110",
"01010011000001000000000000110001",
"00000000001100100000110000001101",
"00000101000110000011111000000100",
"00000000001100011101111100001101",
"01001100000011010101001100000100",
"00111110000001000000000000110010",
"00011101000011010000010100001010",
"01010011000001000000000000110010",
"00000000001100101000000000001101",
"00000100111111000011111000000100",
"00000000001100100101100100001101",
"10111101000011010101001100000100",
"00111110000001000000000000110010",
"10001110000011010000010011101110"
)
,(
"01010011000001000000000000110010",
"00000000001100110001010000001101",
"00000100111000000011111000000100",
"00000000001100101100100100001101",
"01110001000011010101001100000100",
"00111110000001000000000000110011",
"00100000000011010000010011010010",
"01010011000001000000000000110011",
"00000000001100111000000100001101",
"00000100110001000011111000000100",
"00000000001100110111111000001101",
"11010110000011010101001100000100",
"00111110000001000000000000110011",
"10001111000011010000010010110110",
"01010011000001000000000000110011",
"00000000001101000010011000001101",
"00000100101010000011111000000100",
"00000000001101000011001100001101",
"01000001000011010101001100000100",
"00111110000001000000000000110100",
"00111010000011010000010010011010",
"01010011000001000000000000110100",
"00000000001101001011000100001101",
"00000100100011000011111000000100",
"00000000001101000101000000001101",
"11011011000011010101001100000100",
"00111110000001000000000000110100",
"10111111000011010000010001111110",
"01010011000001000000000000110100",
"00000000001101010000110100001101",
"00000100011100000011111000000100",
"00000000001101001110101100001101",
"00110100000011010101001100000100",
"00111110000001000000000000110101",
"00010011000011010000010001100010",
"01010011000001000000000000110101",
"00000000001101010110000100001101",
"00000100010101000011111000000100",
"00000000001101010011101100001101",
"10010110000011010101001100000100",
"00111110000001000000000000110101",
"01110000000011010000010001000110",
"01010011000001000000000000110101",
"00000000001101011101000000001101",
"00000100001110000011111000000100",
"00000000001101011010001000001101",
"00000110000011010101001100000100",
"00111110000001000000000000110110",
"11011100000011010000010000101010",
"01010011000001000000000000110101",
"00000000001101100100001100001101",
"00000100000111000011111000000100",
"00000000001101100100101100001101",
"11111101000011010101001100000100",
"00111110000001000000000000110110",
"01110010000011010000010000001110",
"01010011000001000000000000110110",
"00000000001110000110011000001101",
"00000100000000000011111000000100",
"00000000001101110000110000001101",
"11000101000011010101001100000100",
"00111110000001000000000000111000",
"01110011000011010000001111110010",
"01010011000001000000000000111000",
"00000000001110010010100100001101",
"00000011111001000011111000000100",
"00000000001110001101010100001101",
"01011100000011010101001100000100",
"00111110000001000000000000111001",
"00110100000011010000001111010110",
"01010011000001000000000000111001",
"00000000001110011000111100001101",
"00000011110010000011111000000100",
"00000000001110010110011100001101",
"10000111000011010101001100000100",
"00111110000001000000000000111011",
"10011000000011010000001110111010",
"01010011000001000000000000111001",
"00000000001110111011101100001101",
"00000011101011000011111000000100",
"00000000001110111000101100001101",
"11010001000011010101001100000100",
"00111110000001000000000000111011",
"11011011000011010000001110011110",
"01010011000001000000000000111011",
"00000000001111000100001100001101",
"00000011100100000011111000000100",
"00000000001111001000011000001101",
"00111001000011010101001100000100",
"00111110000001000000000000111101",
"10111011000011010000001110000010",
"01010011000001000000000000111110",
"00000000001111101111110000001101",
"00000011011101000011111000000100",
"00000000001111101110110100001101",
"01100001000011010101001100000100",
"00111110000001000000000000111111",
"00001011000011010000001101100110",
"01010011000001000000000000111111",
"00000000001111111001000100001101",
"00000011010110000011111000000100",
"00000000001111110110101100001101",
"11000010000011010101001100000100",
"00111110000001000000000000111111",
"11110011000011010000001101001010",
"01010011000001000000000000111111",
"00000000010000010001101100001101",
"00000011001111000011111000000100",
"00000000010000000111010000001101",
"01000111000011010101001100000100",
"00111110000001000000000001000001",
"00100001000011010000001100101110",
"01010011000001000000000001000001",
"00000000010000010110010100001101",
"00000011001000000011111000000100",
"00000000010000010100111100001101",
"10010110000011010101001100000100",
"00111110000001000000000001000001",
"01110101000011010000001100010010",
"01010011000001000000000001000001",
"00000000010000011011001000001101",
"00000011000001000011111000000100",
"00000000010000011010010000001101",
"11010001000011010101001100000100",
"00111110000001000000000001000001",
"11000000000011010000001011110110",
"01010011000001000000000001000001",
"00000000010000011110011100001101",
"00000010111010000011111000000100",
"00000000010000011101100100001101",
"00011111000011010101001100000100",
"00111110000001000000000001000010",
"00100110000011010000001011011010",
"01010011000001000000000001000010",
"00000000010000100010101100001101",
"00000010110011000011111000000100",
"00000000010000100010100000001101",
"00111111000011010101001100000100",
"00111110000001000000000001000010",
"00111101000011010000001010111110",
"01010011000001000000000001000010",
"00000000010000100101010000001101",
"00000010101100000011111000000100",
"00000000010000100101001000001101",
"10000111000011010101001100000100",
"00111110000001000000000001000010",
"01100011000011010000001010100010",
"01010011000001000000000001000010",
"00000000010000101010001100001101",
"00000010100101000011111000000100",
"00000000010000101001010100001101",
"11000000000011010101001100000100",
"00111110000001000000000001000010",
"10111000000011010000001010000110",
"01010011000001000000000001000010",
"00000000010000110011100100001101",
"00000010011110000011111000000100",
"00000000001110111011101100001101",
"00000000001111100101011000000100",
"00001010010101000100011000000011",
"01000011100011010000110100000001",
"00111110010101100000010000000000",
"01011000010001100000001011110011",
"01000000010001100000000100001010",
"10001000000011010101010100001000",
"00111110000001000000000001000011",
"10101000010001100000001001010010",
"10000011000011010101010100001010",
"00111110000001000000000001000011",
"01000000010001100000001001000110",
"01111110000011010101010100001001",
"00111110000001000000000001000011",
"01001000010001100000001000111010",
"01111001000011010101010100001001",
"00111110000001000000000001000011",
"01001100010001100000001000101110",
"01110011000011010101010100001001",
"00111110000001000000000001000011",
"01010101010101100000001000100010",
"00000000010000110110100000001101",
"00000010000110000011111000000100",
"00001101010101010000001001011010",
"00000100000000000100001101011110",
"01000110000000100000110100111110",
"00001101010101010000101001011000",
"00000100000000000100001110001101",
"01000110000000100000000100111110",
"00001101010101010000101001010100",
"00000100000000000100001101010111",
"01000110000000011111010100111110",
"00001101010100100000101010010000",
"00000100000000000100001101001110",
"01000110000000011110100100111110",
"00001101010100100000101010001100",
"00000100000000000100001101000110",
"01000110000000011101110100111110",
"00001000000000101111111111010100",
"00000000000000000000110101010110",
"00010100000000000000010000000000",
"01000110001100001110000000111110",
"00001000000000101111111111010100",
"11110000000000001000110111010110",
"10010100100000000000001111111111",
"01000110000001000100000001000110",
"01000110000000010000100101000000",
"01000100010001100000010000000000",
"01000110010101100000000100001001",
"01010110000000010000101010011100",
"00000001000010101010000001000110",
"00001010101001000100011001010110",
"01001100010001100101011000000001",
"01000110010101010000000100001010",
"01010110000000010000101001010000",
"00000001000010010100100001000110",
"00001001010011000100011001010110",
"01011100010001100101011000000001",
"00000000010001100000000100001010",
"00001001010001000100011000000100",
"00000100010000000100011000000001",
"00000001000010010100000001000110",
"11111111110100000100011001010111",
"00000000000100000100011000000001",
"00001001100100001001000101010110",
"11111111110110000100011000001110",
"10111000101011011001100000000001",
"11111111111101001100001010011111",
"00100100111000000000110110001001",
"00111110010010010000010000000000",
"11001110000011010000001100111110",
"01001000000001000000000000100100",
"00001101000000110011010100111110",
"00000100000000000100001011001100",
"00000011001011000011111001000111",
"00000000000011110011000000001101",
"00100011001111100101011000000100",
"11111111110100000100011000000011",
"00011111111111100100011000000010",
"11111111110100000100011000011100",
"00011101000111110011111000000001",
"00001010010010000100011001010110",
"11010100010001100101010100000001",
"11100100001111100000000111111111",
"11000010000011010000100000011011",
"00011110000001000000000000001110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"10010011001111100010001000000100",
"11101110001111100101010100000100",
"11111111110101000100011000100001",
"01001000010001100000100000000010",
"01000110010101100000001000001010",
"01010101000000010000101001001000",
"00000001111111111101010001000110",
"00100001110101110011111001010111",
"00000000111111110100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"11011100010000001111010000101110",
"11111110010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000110001000010",
"00001010100000000100011001010110",
"00100000001011000011111000000001",
"00000000000000001100011001000000",
"00101101000000001111110101000110",
"00000111010000100000101000101100",
"00100011001111100000100000000000",
"00000000101101010100000000101000",
"00000000111111000100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000001000",
"01000000000010000001101101101111",
"01000110000000000000000010100011",
"00101100001011010000000011111011",
"00000000000001110100001000001010",
"00000010101001100011111000001000",
"00000000000000001001001001000000",
"00101101000000001111101001000110",
"00000111010000100000101000101100",
"00011001001111100000100000000000",
"00000000100000010100000000011011",
"00000000111110010100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"01110000010000000011010101111100",
"11111000010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000011101000010",
"01000000001011110100010000111110",
"01000110000000000000000001011111",
"00101100001011010000000011110111",
"00000000000001110100001000001010",
"00101111010001110011111000001000",
"00000000000000000100111001000000",
"00101101000000001111011001000110",
"00000111010000100000101000101100",
"01011010001111100000100000000000",
"00000000001111010100000000101111",
"00000000111101010100011000000000",
"01000010000010100010110000101101",
"00111110000010000000000000000111",
"00101100010000000000000111001000",
"11110100010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000011101000010",
"01000000001000000011011100111110",
"01000110000000000000000000011011",
"00101100001011010000000011110011",
"00000000000100000100001000001010",
"00000000000000000000110100001000",
"10000000010001101000000000000000",
"01100111001111100000000100001010",
"00000000000000010100000000011111",
"11111110111101010100000000001000",
"00000000000000000000000000111101",
"11111111111111111101100010001101",
"11010011100000101000111000000010",
"10001110100101111001101010011010",
"00010000100111010000000100010000",
"10001000000100001001110100000001",
"10001000100000011000111100000001",
"01001101000000000000110000111101",
"01001001010011000100110001001001",
"01001111010000110100010101010011",
"00001001010100110100010001001110",
"01000101010100100101000000000000",
"01001001010100110100100101000011",
"00000000000010010100111001001111",
"01010101010001000100111101001101",
"01001111010101000100010101001100",
"01000100000000000000011101010000",
"01010100010101000100001101001001",
"00000000000001000101000001001111",
"01000101010100110100000101000010",
"01010000010100110000000000000100",
"00000000000001000100111001000001",
"01000101010100100100010101001000",
"00011001000011100001111000001110",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"10010001010101100001111000001010",
"00000100000011110000100110010000",
"00110101000101110000010000001111",
"00001010000000000000010001000010",
"00001000001111011000100100001010",
"00011000000010001001000000011000",
"10101101100110001000100000010000",
"11100101110000101001111110111000",
"01010110000010011000100111111111",
"01100011000000000000011000111101",
"01110100011000010110010101110010",
"00000000000000000000110101100101",
"11011000000011010000001100000000",
"00000010000000101111111111111111",
"01000000000010011001000010010001",
"00010001100100000000000000101000",
"11111111010001100000001000011101",
"00101101000100000001110000000000",
"10001000000100000000101000101100",
"01000010000111000010001000101100",
"00010000000011110000000000001110",
"11111111100111000011111000000010",
"00000000000001000100001000101100",
"00111101100010010001000000001001",
"10010000000110100001101001010011",
"10111000101011011001011000001000",
"11111111110100101100001010011111",
"00010111000011100000100010001001",
"00111110010101100000111000111101",
"01000010001101011111111110110111",
"00110101000010100000000000000010",
"11111111111100010011111000111101",
"01010110000000000000010001000010",
"00001000000000010001110100001111",
"00000000000000000000010000001101",
"00000000000000000000110100000011",
"11011000000011010000001100000000",
"00000010000000101111111111111111",
"00001001100100001001000100011101",
"00010000000000000001000101000000",
"00000000000001100100001000000010",
"01000000100010010001000000001000",
"00011010010100110000000000001101",
"10010110000010001001000000011010",
"11000010100111111011100010101101",
"01010101100010011111111111101001",
"00001101000101110001101000011010",
"00000010111111111111111111011000",
"00000000000001000011110100000001",
"01000100010011100100100101000110",
"10010000000111010000111100110110",
"00000000111111110100011000000010",
"10000010100111010001110000011100",
"00101100001011010101011000000000",
"00000000000001110100001000001010",
"00111101100010000000100000001000",
"00000000000000000011111101000000",
"00001010001011000010110101010011",
"00001000000000000000011001000010",
"00110001010000000011110100001000",
"00101101010100010000000000000000",
"00010100010000100000101000101100",
"11001100100011010000100000000000",
"10000001000000101111111111111111",
"00001101000111010001110100011101",
"00000010111111111111111111011000",
"00010101010000000011110100000001",
"00101101010100000000000000000000",
"00001100010000100000101000101100",
"11111100100011010000100000000000",
"10000001000000101111111111111111",
"00000001010000000011110100001000",
"00010000000010000000100000000000",
"00000000000001100011110110001000",
"01100111011100100110111101100110",
"00111110010101110111010001100101",
"00101100000010100010001001001101",
"00000000000010110100001010010000",
"11110000001111100101000100001110",
"10011100100100000011010111111110",
"00001000111111111000010100111110",
"11000010000000100100011000111110",
"11000010000011010000000000001000",
"01000000000001000000000000001110",
"10111001000011010000000000000101",
"00111110000001000000000000001110",
"00001110000111100000001000110011",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000001101110000011111000100010",
"01000110000000000000011100111101",
"01000101010011000100100101000001",
"00000000000000110011111001000100",
"00000111001111100100101101001111",
"01000101010110000100010100000000",
"01000101010101000101010101000011",
"00011010000110100001110001000111",
"00011100010001110011110100000001",
"00111101000000100001101000011010",
"01000101010100110000000000001001",
"01000011010001010101011001010100",
"00111110010100100100111101010100",
"00001001001111011111110000110101",
"01010100010001010100011100000000",
"01010100010000110100010101010110",
"01001111010001100101001001001111",
"00011110010000100000010000001010",
"11111001001111100100011100000000",
"00000000000101000100011000000000",
"01010110000000010011110000111110",
"01000110001000100111011100111110",
"11101001001111100000000000011001",
"00001010011101000100011000000000",
"11111111111111000000110100000010",
"00111110000000010000001011111111",
"00000100001111011111101111110001",
"01001001010101010101000100000000",
"00000001000011100101101001010100",
"01000001000000000000010100111101",
"01010100010100100100111101000010",
"11111111110101000100011001000011",
"00001111011111010000110100000010",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000001001010000011111000100010",
"11111111111111111110010000001101",
"00010000010001100000001000000010",
"11111111111001000000110100000000",
"00010000000000010000001011111111",
"00001101000101001111010000111110",
"00000010111111111111111111100100",
"11011000010001100000111000000001",
"11010100010001100000000111111111",
"01000000000011010000000111111111",
"01010110000000000000111101000010",
"10011000000010011001000010010001",
"11000010100111111011100010101101",
"01000100100010011111111111111001",
"01110101000000000010001100111101",
"01100110011001010110010001101110",
"01100100011001010110111001101001",
"01110011011011100110100100100000",
"01100011011101010111001001110100",
"01101110011011110110100101110100",
"01100011011011110110110000100000",
"01100100011001010111010001100001",
"01100001011001010110111000100000",
"00000000000001110010000001110010",
"01010100010001100100111101010011",
"01000110010101000100111001001001",
"11000110000000101111111111010100",
"01000100110001100000101001000000",
"00010000000000100001000100001010",
"00000000000110000100011000000010",
"00000010111111111110110001000110",
"00101100000101110001110000001111",
"01000010000111000011100000001111",
"00010111010101000000000000011100",
"00000000010000000100011000001111",
"11100000010001100000011000010110",
"00001010100100010000000111111111",
"01000110000111101000100000010000",
"10010001000111000000001111111111",
"01000000100010000001000000001010",
"00000001000100001111111111010011",
"01000110100010010000000100010001",
"00111101000000011111111111010100",
"00000010000010100100010001000110",
"00010111000001000000000001000110",
"11110011001111100011110100101010",
"11111111111110100100001011111111"
)
,(
"01000110000000000001100001000110",
"00001111000000101111111111101100",
"01000110001011000001011100011100",
"00101100000000100000101001000100",
"00000000000001110100001000011100",
"00000001111111111110000001000110",
"11000110000000000010000001000000",
"11000110100000101111111111010100",
"10000010100011100000101001000100",
"00000010000010100100000001000110",
"11111111010001100001011000010000",
"01000000010001100001110000000011",
"10011110000001010001011000000000",
"11000110100010001000000110001111",
"00111101100000011111111111010100",
"01001101010001010000000000000101",
"01000110001111110101010001001001",
"00001110000111000000000011111111",
"00010111000000000001101101000110",
"00000100010000100001111100111000",
"00000001000000000100011000000000",
"11111111101000100011111000100010",
"10010000100100010101011000111101",
"00000000000001110100000000001001",
"11011110001111100000010000001110",
"10101101100110000001100011111111",
"11110011110000101001111110111000",
"00111101000010001000100111111111",
"00011101010110110011111001010101",
"11111111100000100011111001010110",
"01000110111111111101111000111110",
"01111001001111100000000000011010",
"01001010001111100101011111111111",
"00111110010101010011110100011101",
"00111110010101100001110101000101",
"10110010001111101111111101101100",
"00000000000110100100011011111111",
"01010111111111110110001100111110",
"00111101000111010011010000111110",
"01011001010101000000000000000100",
"00111110010101010100010101010000",
"00111110010101100001110100101001",
"10010001010101101111111101010000",
"00000111010000000000100110010000",
"00000000001000000100011000000000",
"10011000111111111000110000111110",
"11000010100111111011100010101101",
"01000110100010011111111111110011",
"00110101001111100000000000011010",
"00000110001111100101011111111111",
"00000000000001000011110100011101",
"01010100010010010100110101000101",
"11111111110011100011111001010101",
"01010011000000000000011000111101",
"01000101010000110100000101010000",
"11101110001111100101010101010011",
"00010101001111100101011000011100",
"01011010001111100100100111111111",
"01010110001111100100110011111111",
"00000000000110100100011011111111",
"01010111111111110000011100111110",
"00111101000111001101100000111110",
"01010000010100110000000000000101",
"01010101010001010100001101000001",
"01010110000111001100110000111110",
"00111110001001000000110000111110",
"00111110010101111111111101100110",
"00111110010101110010010000000101",
"00000010001111010001110010111101",
"01010011010100100100001100000000",
"01010011000010110101001100001011",
"00111110000010110101001100001011",
"10010000100100010000000000011001",
"10010001000001000001001100111110",
"10010001000100000001011100001010",
"10001001000100000010011000001010",
"00111101100010010001000000010001",
"01010010010100000000000000000101",
"11000110010101000100111001001001",
"00001111100000101111111111010100",
"01011100000101110101010100001111",
"00000001000001100100001000100010",
"11000110101101101001000111010101",
"00010000100111000000000000100000",
"00001111000000000000011101000010",
"01000000000101110011011000001111",
"10010110000011100000000000000001",
"10011100100110011000111010010000",
"00010000110001101001011010101100",
"00001111000011110101011000000000",
"00010110000100000000111101010101",
"01011011000101110000101000100000",
"00000000000000100100001000011111",
"10101011100110110001011000010000",
"10001000111111111110101111000010",
"01000110000010011001011010010000",
"00010111000100000000000001000000",
"00001111000000110001011000111110",
"10001111010000100010001000001111",
"00001101000011110000111100000000",
"01111111111111111111111111111111",
"00010111000010101001000101010111",
"00100110000010101001000100010000",
"10010000001000011000100100010000",
"00100110000011110101011000001000",
"01010001100010000001000000001010",
"00001001100100001001000101010110",
"01010011011000010000111100001111",
"01100001000010110101001100001011",
"01100010011000100110001001100010",
"00001000100100000010000100001001",
"00001010001001100000111101010110",
"01100001011000011000100000010000",
"01100010011000100110001001100010",
"10010001000011110000111100001001",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"10011111101110001010110110011000",
"10001001111111111101000111000010",
"00001010100100010000111100001111",
"00001010100100010001000000010110",
"01010110100010010001000000100101",
"00010111000010101001000101010011",
"00100110000010101001000100010000",
"00001111000011111000100100010000",
"01010011000010110101001101100001",
"01100010011000100110000100001011",
"01010001000010010110001001100010",
"10010001000010110101000100001011",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"01000010000111110010101000001111",
"10010000000010011111111111010111",
"00010000000010100000101000001000",
"00000000000000010100000010001000",
"00001111000011110110000100011000",
"01100010011000100110001001100001",
"10010000100100010000100101100010",
"00010000000101110000101010010001",
"00010000001001100000101010010001",
"01010101000010001001000010001001",
"01010101100010000001000000100011",
"10001001000100000001000100101000",
"00010000000101100000101010010001",
"00010000001001010000101010010001",
"00011001100010000001000010001001",
"01000000000000101010000100111110",
"00101100000010100000000000001010",
"00001001000000000000010101000010",
"01010111001000110101010101010111",
"10000001111111111101010011000110",
"01010101000000000000011100111101",
"01001101010001000010111101000100",
"00001110100100000100010001001111",
"00111110100010000001000000010111",
"10010000100100011111111010101001",
"00010000000100010000101000001001",
"11101101001111100011110110001001",
"00000110001111010000101011111111",
"00101111010001000101010100000000",
"10010000010001000100111101001101",
"00101010000011111001000100001000",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00000001010000100010100100010001",
"11011001001111100010000100000000",
"11000010101010101010010011111111",
"10010000001000010000000000000110",
"10001000000100000010000100001000",
"01010101000000000000011000111101",
"01001111010011010010111101001101",
"11001110001111101001000001000100",
"00101001000010001001000011111111",
"00010001000000000000100101000010",
"00000000000000010100001000101010",
"10011001000101100001000100100001",
"00000110001111011000100100010000",
"00101111010011010101001100000000",
"10010001010011010100010101010010",
"01000010001010011010010010010000",
"10010001001000010000000000000001",
"00101001100010000001000000001010",
"00100001000000000000000101000010",
"10101010000000000001011000111110",
"00100001000000000000100111000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"01000110000000000000011000111101",
"01001111010011010010111101001101",
"11111111110101001100011001000100",
"01100001000011110101011010000010",
"01100001000011110101011000001000",
"00001001011000100110001000001000",
"11010100110001100110001001100010",
"00000010001111011000000111111111",
"00111110001010100100110100000000",
"00111101000010101111111110111001",
"00101010100100000000100010010000",
"10001000000100001000100000010000",
"00111101111111110110000000111110",
"00111110001010100000000000000001",
"00111101000010101111111111101110",
"01001101001011110000000000000100",
"11100011001111100100010001001111",
"00000001001111010000100011111111",
"00001000100100000010111100000000",
"00010000111111111001000000111110",
"11111111001111110011111010001000",
"01001101000000000000001100111101",
"11101101001111100100010001001111",
"00000101001111010000101011111111",
"01001101001011110010101000000000",
"00000100000011110100010001001111",
"00101101000000000010110101000110",
"00000101010000100000101000101100",
"01000000100011101101011100000000",
"10010000110101100000000000000111",
"10010111000000000010101111000110",
"00000110110000100000100010101100",
"00001000100100000001100100000000",
"10010000100010000001000000011000",
"10010011110000101011011100001000",
"01000110000001001001000000000000",
"00101010001011010000000000110000",
"00111001010001100000111100001010",
"00100010001110000001011100000000",
"00000000001100000100011000011111",
"01000001010001100001011100011100",
"00001010001010100010110100000000",
"00000000010110100100011000001111",
"00011111001000100011100000010111",
"00011100000000000011011101000110",
"00000000011000010100011000010111",
"00001111000010100010101000101101",
"00010111000000000111101001000110",
"01000110000111110010001000111000",
"00010111000111000000000001010111",
"11111111111111111110010000001101",
"00101010001011010000001000000010",
"00000000000001100100001000011111",
"01000000100010000001000000001001",
"10010000100100010000000001000110",
"00001001100100001001000100001001",
"00010000000100010000111001010110",
"00100011110000101011010110001001",
"00001110000011101001101100000000",
"00000000000011100100001000100110",
"00001010100100011001000010010001",
"00001010100100010001000000010110",
"00010001100010010001000000100101",
"00001111000011111000100100010000",
"00010000000101100000101010010001",
"00010000001001010000101010010001",
"11111111110110010100000010001001",
"10001001000100010001000000001001",
"00010000000101100000101010010001",
"00010000001001010000101010010001",
"00011000100010000001000010001001",
"11111111011010010100000010011001",
"00001010100100011000101000010001",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00111101100010010001000100010000",
"00101111001010100000000000000010",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"00111101000010001111111100100000",
"01001110001111100000000000000111",
"01000101010000100100110101010101",
"00000111010000100010100101010010",
"01010100001111100010000100000000",
"00000000010001110100000000000000",
"00101101000000000100000001000110",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"10010001000010001001000000001000",
"01000110100010100001000110101010",
"00111000001011010000000000011111",
"00010111000000000000111001000010",
"00010001000010011001000000011001",
"10001000000100000000101010010001",
"11101010010000001000100000010000",
"00100011100100000000100011111111",
"00000000001000000100011000001111",
"00100010001000000001011100010000",
"10001000000100000000101010010001",
"01000110000100010010001100010000",
"10001001000100000000000000100000",
"10010001001000100010000000010111",
"00111101100010000001000000001010",
"01001111010000110000000000000111",
"01010010010001010101011001001110",
"00000111010000100010100101010100",
"10011100001111100010000100000000",
"00000000001110110100000011111111",
"00101101000000000100000001000110",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"00000000000111110100011000001000",
"00001111010000100011100000101101",
"10010000000110010001011100000000",
"00010000000010101001000100001000",
"00010000000101110000111010001000",
"11111111111010010100000010001000",
"00100000100100011001000000001000",
"10001000000100000000101010010001",
"01000110000100000010000000010001",
"00010111000100010000000000100000",
"00001010100100010010001000100011",
"00111101100010011000100000010000",
"01010011010000010000000000000110",
"01010100010001100100100101001000",
"00000000000001110100001000101001",
"11111111101010010011111000100001",
"01000110000000000011101001000000",
"00111000001011010000000001000000",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"00101101000000000001111101000110",
"00000000000011110100001000111000",
"00001000100100000001100100010111",
"00001010100100010001011100001110",
"10001000000100001000100000010000",
"00001000111111111110100101000000",
"01000110000011110010001110010000",
"00010111000100000000000000100000",
"00001010100100010010001000100000",
"10001000000100001000100000010000",
"00010000000010101001000100100011",
"00000000000001100011110110001000",
"01000110010010010100100001010011",
"11010100110001100100110001010100",
"00001111100100011000001011111111",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00001111100100010110000110001000",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"10101010101001000110000110001000",
"01100010000010010110001001100010",
"00000000000010011100001001100010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"11111111110101001100011010001000",
"00000000000001100011110110000001",
"01000110010010010100100001010011",
"00001111100100010101001001010100",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00001001100100011001000010001000",
"01000010001010100000111110010001",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"00010001100010000001000000001010",
"10100100100010100001000110001010",
"10101010111110110111000000111110",
"00100001000000000000100111000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"00001010000010100000100010010000",
"00000010001111011000100000010000",
"10010001001010100100010000000000",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10010001100100001000100000010000",
"00101010000011111001000100001001",
"00100001000000000000100101000010",
"00001111010101100000100010010000",
"10001000000100000000101000100110",
"10001010000100011000101000010001",
"11111011001011110011111010100100",
"00001001110000101010101000001001",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"00000010001111011000100000010000",
"10010000001011110100010000000000",
"00000000000000000000110100001000",
"00010000001001001000000000000000",
"00000000000001000011110110001000",
"01000100010011110100110101000100",
"00101100001000100000111100001111",
"00111101000000000000000101000010",
"00001111010000100010101000001111",
"00001100001111111100011000000000",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00000000000000110100000010001000",
"10011001000001000011111111000110",
"00001010100100010000111100001111",
"00001010100100010001000000010110",
"01000011100010010001000000100101",
"01001010111111111111000001000010",
"00010100010001100000111100100011",
"10010000001000100010000000000000",
"00010001001000110100101000001000",
"00100000000000000001010001000110",
"00111101100010010001000000100010",
"01001110010001100000000000000111",
"01010100010000010100011101000101",
"10010001000010001001000001000101",
"00000000000011010000100110010000",
"01010110001111111111000000000000",
"10001000000100001000101111010100",
"00000000000000010100001000101001",
"00100010010000100000111000100001",
"01000010010000110001101100000000",
"10010001000100010000000000001001",
"11110000001111100001000100001010",
"00010001100010000001000000000000",
"00010001000010101001000110001010",
"00111110000011110000111110001010",
"00001010100100010000000011100011",
"00001010100100011000101000010001",
"00001000111111111101101001000000",
"00001111110000101010101010001001",
"00001001100100001001000100000000",
"11110000000000000000000000001101",
"00010000000100010101011000111111",
"00000011000010100011111010001001",
"01000100000000000000001100111101",
"10010001100100000100011000111110",
"00010000000011100101011000001001",
"10011101001111101000100100010001",
"00000100000011111001000011111100",
"00010111000000000010111001000110",
"00011100001101100000111100101100",
"10001000000000000011001001000010",
"00011000000010001001000000011001",
"00001111100100010000100010010000",
"00000000000010010100001000101010",
"01010110000010001001000000100001",
"00010000000010100010011000001111",
"00010001100010100001000110001000",
"10010000111111000111001100111110",
"10010001100010100001000100001000",
"00001001010000100010101000001010",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"00010001000100001000100000010000",
"10100001100101111001000010001001",
"00111110000010011001000110010000",
"00000100000100001111111100001010",
"00101101000000000100010101000110",
"01000110000011110000101000101100",
"00101100000101110000000001100101",
"00110110000100010000101000100010",
"00000000000100000100001000011100",
"00011000000100000000111001010110",
"00111110100010010001100100010001",
"10010000000010011111110000110100",
"00001001100100011001000010010110",
"11100100000011010101011010001001",
"00000010000000101111111111111111",
"00010000111111101101100100111110",
"11111111001000010011111010001000",
"01010111000000000011001000111110",
"01100010011000010110000100111101",
"10010001011000100110001001100010",
"01001011000010001001000000001001",
"00010101010001100001000000100000",
"00010000001000100010001100000000",
"00010001010101100010000001001011",
"00000000000101010100011010001001",
"10010001001001010101011000100011",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00111110000000000000011000111101",
"01000001010011110100110001000110",
"11111111110101001100011001010100",
"10010000000010001001000010000010",
"00001111111111111111111110001101",
"00000000000011011001110000000000",
"00011100111111111111000000000000",
"00000000000000000000110100001110",
"00110110000111000111111111110000",
"10001101000000000000011001000010",
"00000000000100000000000000000000",
"10010001000010101001000110100010",
"11111111100011010001000000001010",
"10011100000000000000111111111111",
"11110000000000000000000000001101",
"00001101000011100001110011111111",
"01111111111100000000000000000000",
"00000110010000100011011000011100",
"00000000000000001000110100000000",
"10010000101000100000000000010000",
"00000000100011011010010010010001",
"10011100100000000000000000000000",
"11110000000000000000000000001101",
"10010001000110110001110001111111",
"00001101100010000001000000001010",
"01111111111100000000000000000000",
"00001101000101100001101100011100",
"00011111111110000000000000000000",
"00000000000000000000110100010111",
"00111000001011010011111111110000",
"00000000000100100100001000001010",
"00000000000011011001101000001000",
"01010101111111111110000000000000",
"10001001100010000101011000101000",
"11111111110101001100011010001001",
"00101101010101100011110110000001",
"00000000000001000100001000101010",
"10001000000100000000101010010001",
"00001000100100000001101000001000"
)
,(
"00010001100010100001000110100010",
"10010001000011110000111110001010",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"10001010000100011000101000010001",
"00001111111111110010011000111110",
"00010000000000000000000000001101",
"00001010001010100010110100000000",
"10001101000000000000011001000010",
"10000000000000000000000000000000",
"11111111111111110000110110011100",
"00111000000101110000000000011111",
"10010000000000000000110101000010",
"10101000110101010001101100001000",
"00000000100011011000100000010000",
"10010110000000000001000000000000",
"11111111000011010000100010010000",
"00011100000000000000111111111111",
"10001001000100000010001000010001",
"10000001111111111101010011000110",
"00001000100100001001000100111101",
"00001111111111111111111100001101",
"00001101000100010001110000000000",
"01111111111100000000000000000000",
"00000110010000101001000000011100",
"00000000000000000000110100000000",
"00010001001000100000000000010000",
"00001000100100000001101010001010",
"10001000000100000010010100001110",
"00001001010000100010101000010001",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"10001001000100001000100000010000",
"01000110000000000000001000111101",
"00000000001100100100011000101010",
"00001000100100000010101000010111",
"00010000000100010000101010010001",
"00010101010001100001101010001001",
"00001000100100000010001100000000",
"00010000000100010000101010010001",
"00010101010001100001101010001001",
"00001111000011110010001100000000",
"00000001010000100010100100010111",
"00110110010001100010000100000000",
"00001111001010100001011100000000",
"00001010000010100001110000110110",
"10010000100100010011110100011100",
"11111111100100010011111000001001",
"00001010100100011000101000010001",
"10001000001111101000101000010001",
"00010001000010001001000011111111",
"00100011000000000001010001000110",
"00000000000101000100011000010000",
"01000010001010010001011100100011",
"10010001100010100000000000001111",
"00100001000010101001000100001010",
"00010000111110110101111000111110",
"00000100010000001000100100010001",
"01010100001111101000100000000000",
"00010110000010101001000111111011",
"00100101000010101001000100010000",
"00001111100110101000100100010000",
"00001000101010001101010100011010",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"00001111000011111000100000010000",
"00000110010000100010110000100010",
"00000000000000001000110100000000",
"00001111100111001000000000000000",
"00100000000000000000000000001101",
"00010000001010100001011100000000",
"00010100010000100001110000011010",
"10010001000011110000111100000000",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"00010000000000000000000010001101",
"11011110010000001001011100000000",
"01010100100010000001000011111111",
"00001001100100001001000101010110",
"00001101000011110000100010010000",
"00000000001111111111111111111111",
"00011010000100000011100000010111",
"11100000000000000000000000001101",
"00011100001101100001011111111111",
"10010000000000000000110101000010",
"10001000000100000001101100001000",
"00000000100011010010100001010101",
"10010110000000000001000000000000",
"10010001000110000000111001010110",
"10010001000100000001011000001010",
"10001001000100000010010100001010",
"10001000000100000001110001011000",
"10011111101110001010110110011000",
"10001001111111111100010111000010",
"00001000100100000000100010010000",
"01010101100010000001000000011011",
"11111111000011010000111100101000",
"00010111000000000000111111111111",
"00101100000110100001000000111000",
"00000000000001100100001000011100",
"00010000000000000000000010001101",
"00001000100100001001011000000000",
"00001111111111111111111100001101",
"00100010000100010001110000000000",
"00111110001111011000100100010000",
"00001101001111101111110001010001",
"00000000000000100011110111111111",
"00001000001111100010101101000110",
"11111101101101010011111000000000",
"01000110000000000000001000111101",
"00001001100100001001000100101101",
"00000000000011010001000101010110",
"00011100100000000000000000000000",
"00010101010001100001101000010001",
"11111111010001100010001100000000",
"01000110000111110001011100000011",
"01000110000101100000001111111110",
"01010101001000000000000000010101",
"11010110100100000010001000100011",
"01010010000100010000111101010110",
"11111110101000010011111000001011",
"00010101010001100001101000010001",
"11111111010001100010001100000000",
"00011100001010100001011100000111",
"00010001000000000010001001000010",
"10111101001111101000100100010000",
"00001111000011110000111111111110",
"00111110000011110000111100001111",
"00010000000100011111110101100111",
"00111110111111010110001000111110",
"10010000100100011111111110011001",
"00011000000010110101010000001001",
"11001000010000000000110001010100",
"10010001000010001001000011111111",
"10001001000100000001000100001010",
"00111101100010011000100100001000",
"00101111010001100000000000000010",
"00000000000000000000110100001111",
"00001101000111001000000000000000",
"00111111111000000000000000000000",
"10000001001111100101011000100010",
"00000000011111010011111011111110",
"00001111000000000000000000000000",
"11110000000000000000000000001101",
"00010100010001100001110001111111",
"11111111010001100010001100000000",
"01000010001010010001011100000011",
"00001001000010000000000000000111",
"01010011010000000000111001010110",
"00000000001111100100011000000000",
"01000010000010100011100000101101",
"00101010000010010000000000010111",
"00001101000000000000100101000010",
"10000000000000000000000000000000",
"00000000000001100100000001010110",
"11111111111111111111111100001101",
"00110011010000000101011101111111",
"00001001100100011001000000000000",
"11111111111111110000110110010000",
"00001101000111000000000000001111",
"00000000000100000000000000000000",
"00010001100010100001000100100010",
"00010111000000000011010001000110",
"00000000000001100100001000110111",
"01000000111110100000011000111110",
"00111110001000010000000000000100",
"11000010101010101111101001001110",
"10010000001000010000000000001001",
"00100110000011110101011000001000",
"10001000100010000001000000001010",
"01010010000000000000101000111101",
"01010000010010010100001101000101",
"01000001010000110100111101010010",
"00000000000011010000111101001100",
"00011100011111111111000000000000",
"11110000000000000000000000001101",
"01000010001010010001011100111111",
"00001101000010010000000000001001",
"10000000000000000000000000000000",
"01000110001111010101011000011100",
"11000110001000110000000000010100",
"00001000100100000000000000110100",
"00011000110000101011011110010111",
"00100000110001100101011100000000",
"11000010101010011001011100000000",
"00100000010001100000000000001010",
"00100000000101100001000000000000",
"00000000000001010100000000011100",
"00011100001000000001000000001010",
"00000011001111011000100001010110",
"01000100001111100100011000000000",
"10110100001111100000111100001111",
"10010000100100001001000111111111",
"00100100000010101001000100001000",
"00100010100010000001000010100100",
"00101010000100010001111100101100",
"10010001100010100001000100011100",
"11000010100010100001000100001010",
"00000000000011010000000000001001",
"01010110001111111111000000000000",
"00111101111111101000000000111110",
"01110100011100110000000000000110",
"01100110011100000110100101110010",
"00001011010100010000111100001111",
"01101110001111100000101101010001",
"00100010000110100000111111111110",
"00011100001010100000111100110110",
"00001001010000100001111100001010",
"00001001100100001001000100000000",
"10001001000100000001000100001001",
"00111101000010010000111100001111",
"01001100010001100000000000000101",
"00001111010100100100111101001111",
"01010001000010110101000100001111",
"11111110010001110011111000001011",
"00110110001000100001101000001111",
"00001010000111000010101000001111",
"10010001000000000000100101000010",
"00010001000010010000100110010000",
"00001111000011111000100100010000",
"00000000000001000011110100001001",
"01011000010000010100110101000110",
"00111000001111100000111100001111",
"10010000100100001001000111111111",
"00100100000010101001000100001000",
"00100010100010000001000010100100",
"00101010000100010001111100101100",
"10001010000100010001110000011111",
"10001010000100010000101010010001",
"00001101000000000000100111000010",
"00111111111100000000000000000000",
"11111101000101100011111001010110",
"01000110000000000000010000111101",
"10010001010011100100100101001101",
"00101110001111100000100110010000",
"10001001000100000001000100000010",
"00111110111110111011011000111110",
"00000110001111010000000111001000",
"01001111010100100100011000000000",
"00111110010001000100111001010101",
"11111011000011010000000001010000",
"00001101001111111111100100100001",
"01010100010001000010110100011000",
"00111110111111011101010000111110",
"00000011001111011111101000100101",
"00101010001010100100011000000000",
"00001111000011110000111100001111",
"00001101111110111000101000111110",
"00111111111100000000000000000000",
"11111101101110110011111001010110",
"00111110000000110101101000111110",
"11101010001111101111110011001000",
"00000000000001010011110100000001",
"01001111010000110100000101000110",
"01101011101100010000110101010011",
"00010111000011010100000000000010",
"00111110101110111011010101010101",
"01110101001111101111101101100011",
"00000000000001100011110100000001",
"01001111010000110100000101000110",
"10010000100100010100100001010011",
"11110000000000000000000000001101",
"00010000000100010101011000111111",
"00111110000011110000111110001001",
"01111110001111101111101101000111",
"00000011000111010011111011111101",
"00111110111111011000001100111110",
"00000101001111010000000000101001",
"01001100010000010100011000000000",
"00001111000011110100011101001111",
"00101100001111100000111100001111",
"00000000000000000000110111111011",
"00111110010101100011111111110000",
"11111100001111101111110001110000",
"11111100011010100011111000000010",
"00111101000000011000110000111110",
"01000001010001100000000000000101",
"00001111010011100100100101010011",
"00111110000011110000111100001111",
"10010110001111101111101100001011",
"00001001100100001001000111111001",
"01010110000010011001000010010001",
"00010001000011110001000000010001",
"00010100001111100000101101010010",
"00000000001000100100001011111100",
"00010001100010010001000000010001",
"11111010111011010011111000010000",
"00001011010100101001000010010001",
"00001100010100010000111000011000",
"00101010100100000001100000011010",
"01111011001111101000100000010000",
"11111101000111100011111011111001",
"01000000111111000010001100111110",
"00001000100100001111111111010100",
"00010000000100010000101010010001",
"10001001100010010000100010001001",
"01000110000000000000011000111101",
"01001110010010010101001101000001",
"10010000000010110101001101001000",
"11111101001111101001000100001000",
"11111111101000110011111011111100",
"00000000000101111100001010101010",
"00001001001000011111101100001101",
"00101101000110000000110101000000",
"11000010101010010101010001000100",
"11011010001111100000000000000110",
"00000000000000110100000011111100",
"10001000111110111110011100111110",
"01000110000000000000010100111101",
"01001110010000010101010001000001",
"11110000000000000000000000001101",
"11010101001111100101011000111111",
"00001101000011110000111111111011",
"01000000000000000000000000000000",
"11111100101101110011111001010110",
"00111110111110010000100000111110",
"11100110001111101111110010111100",
"00000000000000000000110100000000",
"00111110010101100011111111100000",
"00000110001111011111101001101011",
"01010100010000010100011000000000",
"00001111001100100100111001000001",
"11111010010111010011111000001111",
"10010001111110001110100000111110",
"00001101010101100000100110010000",
"00111111111100000000000000000000",
"00001111100100001001000101010110",
"00111110000010110101001000010001",
"00100010010000101111101101100011",
"10001001000100000001000100000000",
"00111100001111100001000000010001",
"00011000000010110101001011111010",
"00011010000011000101000100001110",
"10010010001111100001100100001110",
"11111000110011000011111011110101",
"10010001111111000110111100111110",
"11111011011100100011111010010000",
"10010000111111111101010001000000",
"00010001000010101001000100001000",
"10001001000010001000100100010000",
"00000000000001100011110110001001",
"01000001010101000100000101000110",
"00100001001111100100100001001110",
"00001101100100001001000100000000",
"00111111111100000000000000000000",
"10001001000100000001000101010110",
"00111110111111000100001100111110",
"00000000000011011111101101001000",
"01010110001111111110000000000000",
"00111101111110011111001000111110",
"01000011010001100000000000000100",
"10010000100100010101001101001111",
"01010101000010011001000010010001",
"11110000000000000000000000001101",
"00010000000100010101011000111111",
"00001111111110110010011100111110",
"00111110000010110101001000010001",
"00011101010000101111101011101111",
"10001001000100000001000100000000",
"11001000001111100001000000010001",
"00001011010100010101011011111001",
"00001100010100000000111000011000",
"00111110111110000101110100111110",
"10010000100100011111110000000000",
"01000000111110110000001100111110",
"00001000100100001111111111011001",
"00010000000100010000101010010001",
"10001001100010010000100010001001",
"01000110000000000000010100111101",
"01001000010100110100111101000011",
"00001101111111111011001100111110",
"00111111111100000000000000000000",
"11111011110011110011111001010110",
"01000110000000000000010000111101",
"00001111010100000101100001000101",
"00000000000000000000110100001110",
"00101100000111000111111111110000",
"00001010001000100010101000001111",
"00001000000000000000110001000010",
"00000000000011010000100000011010",
"01010101111111111110000000000000",
"10010001001111010101011000101000",
"01000110000110100000100010010000",
"01000110001000110000000000010101",
"10010000000101110000001111111111",
"00111110100010000001000000101010",
"01000010000011011111011111111110",
"00001101001111111110011000101110",
"11111110111110100011100111101111",
"00010001111110010101001000111110",
"00100011000000000001010001000110",
"00010111000001111111111101000110",
"00000000000010010100001000101100",
"11110000000000000000000000001101",
"00001101010000000101011000111111",
"00010001000100000001000100000000",
"11110000000000000000000000001101",
"00111110010101100001110001111111",
"10010001100010011111101101110100",
"00000000000000000000110110010000",
"00111110010101100011111111110000",
"00010000000100011111101101011101",
"11111011011000100011111010001001",
"10001111000010011001000010010001",
"00010000000100010101010110001111",
"00001011010100100001000100001111",
"01000010111110100010101000111110",
"00010000000100010000000000100000",
"00111110000100000001000110001001",
"10010000100100011111100100000011",
"00001110000110000000101101010010",
"00101010100100000000110001010001",
"10010011001111101000100000010000",
"11111011001101100011111011110111",
"01000000111110100011101100111110",
"00001000100100001111111111010110",
"00010000000100010000101010010001",
"10001001100010010000100010001001",
"00111101111110100010101100111110",
"01000101010001100000000000000110",
"00110001010011010101000001011000",
"11110000000000000000000000001101",
"00011001001111100101011000111111",
"11111111001110110011111011111010",
"01000110000000000000001100111101",
"00110010001111100100111001001100",
"01101011101100010000110111111111",
"00010111000011010100000000000010",
"00111110101110111011010101010101",
"00000101001111011111101011111000",
"01001110010011000100011000000000",
"00001111000011110011000101010000",
"10100100001111100000111100001111",
"11110111001011110011111011111000",
"10010001000010011001000010010001",
"00010001010101100000100110010000",
"01010010000100010000111100010000",
"11111001101011010011111000001011",
"00010001000000000010001001000010",
"00010000000100011000100100010000",
"01010010111110001000011000111110",
"01010001000011100001100000001011",
"00011000000011100001101000001100",
"00111110111100111101110000111110",
"10111001001111101111011100010110",
"00111110100100001001000111111010",
"11010100010000001111100110111100",
"10010001000010001001000011111111",
"10001001000100000001000100001010",
"00111101100010011000100100001000",
"01001100010001100000000000000100",
"01101101001111100100011101001111",
"00001101100100001001000111111110",
"00111111111100000000000000000000",
"10001001000100000001000101010110",
"00111110111110101000111100111110",
"00000000000011011111101010000001",
"01010110010000000000000000000000",
"00111101111110101000001100111110",
"01010011010001100000000000000100",
"10010000100100010100111001001001",
"00010001111111111000011100111110",
"11001010001111101000100100010000",
"00000000000001010011110111111101",
"01001110010010010101001101000110",
"00001101000010001001000001001000",
"01111111111111111111111111111111",
"10010001100010000001000000011100",
"00010001010101100000100110010000",
"00000000000000000000110100010000",
"00111110010101100100000000000000",
"00001111000011111111101001010000",
"00000100001111100000111100001111",
"00111110000100000001000111111000",
"00001011010100111111101000111001",
"00000000000011010000101101010011",
"01010110010000000000000000000000",
"00111110111101111111001000111110",
"00111110100100011111101000110100",
"00010000000011111111101000100101",
"00011000000010110101001010001000",
"00111110000011000101000100001110",
"01000010000111111111100011111011",
"00001000100100001111111111010000",
"00010000000100010000101010010001",
"00111101100010010000100010001001",
"01010011010001100000000000000111",
"01001111010000110100111001001001",
"11111111100011100011111001010011",
"00111101111110100000011100111110",
"01010011010001100000000000000101",
"00111110010101000101001001010001",
"10010000100100011111110111001100",
"11110000000000000000000000001101",
"00010000000100010101011000111111",
"10010001111110011110111100111110",
"11111001110111110011111010010000",
"00010001100010010001000000010001",
"11101001001111101000100100010000",
"11111001110111100011111011111000",
"01000110000000000000010000111101",
"10010001010011100100000101010100",
"11000110001111100000100110010000",
"00001101000010001001000011111001",
"01111111111111111111111111111111",
"00001111100010000001000000011100",
"00010001001011000010001000001111",
"00010001000010101001000110001010",
"00001111111110011011000000111110",
"00001111001101100010001000011010",
"00010000000010100001110000101010"
)
,(
"00000101001111010010001010001001",
"01000001010101000100011000000000",
"01001001001111100100100001001110",
"01000010001010010000111000000010",
"00001101001000010000000000000001",
"00000010111111111111111111000000",
"01000010001110000001011100000010",
"00101110010001100000000000010000",
"10000100001111100101010100000000",
"00000001000011010011111000000001",
"01000000000000011011110000111110",
"01000010001010010000000000101101",
"01000000110001100000000000011101",
"00100001100001101000111000001000",
"00001001100100001001000101010110",
"01010110000000000011000001000110",
"10011000000000010110011000111110",
"11000010100111111011100010101101",
"10001111100010011111111111110010",
"01000110010101101000100010000101",
"00011000000011110000000000101110",
"00001000000000010101001000111110",
"01000110000000001101101000111110",
"00001110000111100000100001000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00000000000000100011110100100010",
"10011001001111100111111001000110",
"11101111111111000011111011111111",
"01000110000000000000001100111101",
"11011001001111100010111000101110",
"00000000101101010011111000000001",
"01000110000000001101110000111110",
"00111110010101010000000000101110",
"01011010001111100000000100011111",
"00001000010000000100011000000001",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111101001000100000010000011001",
"00101110010001100000000000000010",
"00111110111111111101011100111110",
"00000100001111011110111111001010",
"00101110010100110100011000000000",
"00000001101001100011111000101110",
"00111110000000001000001000111110",
"10010000000011100000000010101001",
"01010011100010000001000000101010",
"00001000111100011111001000111110",
"00101110010001100001011110010000",
"00011000100010000001000000000000",
"00111110000000001101111000111110",
"01000000010001100000000100011001",
"00011001000011100001111000001000",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"01000110000000000000001100111101",
"11001000001111100010111001010011",
"11101111100010000011111011111111",
"01000110000000000000010000111101",
"00001101001011100010111001000101",
"00000010111111111111111111000000",
"00101101000000000100000001000110",
"00000000000001000100001000111000",
"10001000000100000000101010010001",
"00101010001011010101001100001000",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"00000000000000110011110100000001",
"01000110001011100100010101000110",
"00011000000001100000100001000000",
"01000000010001100001100010010000",
"00010000000000110001011000001000",
"00001000010000000100011010001000",
"00000000000011010011110100000101",
"00101101010101000100010101010011",
"01000011010001010101001001010000",
"01001111010010010101001101001001",
"00001000010000001100011001001110",
"00011001000011100001111000010000",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00011001000101100000111100001111",
"00000000001100000100011000000100",
"01010101000011110010110000010111",
"01000010000111000011100000010111",
"01000000000110010000000000000100",
"00000101000100001111111111101010",
"11000110001111011000100000001000",
"00001000100100000000100001000000",
"00011001000011100001111000010001",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00110000010001100000010000001111",
"00001111001011000001011100000000",
"00011100001110000001011101010101",
"10011001000000000010010001000010",
"00011000000011111001000000011001",
"10001000000100000001100100001110",
"00001001100100001001000101010110",
"00001111000000000000100101000000",
"00001111000001000001011000010000",
"10011000000000110001011000010000",
"11000010100111111011100010101101",
"00001001100010011111111111110001",
"00010001111111111100110101000000",
"10001001000100000000100000000101",
"00001000010000001100011000111101",
"10000100100110011000111010011110",
"10011001100011111010000011001110",
"00010001101000101000010010011001",
"00000000001011010100011000000100",
"00010001000101110010110000010111",
"10010110100011111000111100010110",
"00010000000100010000100010010000",
"00001001100100001001000110001000",
"00010000000000000000011101000000",
"00010000000000111000010010001110",
"10111000101011011001100010001000",
"11111111111100111100001010011111",
"10001000000000110001000010001001",
"10011001100110011000111110011000",
"01000110001111011000100010000101",
"00100110001111100000000001000101",
"00000111010000100010100111111111",
"00101101010001100010000100000000",
"00000000000000110100000000000000",
"00111110000000000010101101000110",
"00000001001111101111111100010101",
"11100100000011010011110100000000",
"00000010000000101111111111111111",
"00110101111100010000110100111110",
"00111110000000000000011001000010",
"00000001010000001111111111110000",
"00000001001111100000100000000000",
"00101101010011010011110100000000",
"00000110010000100000101000111000",
"00000000010101110100011000000000",
"00101001000000000000100001000000",
"00100001000000000000000101000010",
"00010110000000000011000001000110",
"00111101111111101110000000111110",
"01111001001111101001000110010000",
"00111110000011110000111111110111",
"00001111000011111111100001111011",
"00001010111101111110010100111110",
"01011110001111100000100010010000",
"00010001100010100001000111110111",
"11110101000111010011111010010001",
"00010000000100011000100000010000",
"01000110010101100011110110001001",
"00001111000001010000100001000000",
"00000000000010010100001000101010",
"00111110000000000010110101000110",
"10010010001111101111111010101101",
"00000000000011010000111111110011",
"00011100011111111111000000000000",
"00001111000000000000100001000010",
"11111011011001110011111000001111",
"01010110000000000000001001000000",
"11111111111001000000110100001110",
"10010000000000100000001011111111",
"00111110100010000001000000101010",
"10010000100100011111001110000010",
"00111110111110110101000000111110",
"10010011001111101111011100100000",
"10010001000100010000101011110111",
"00001101000100000001000100001010",
"00000010111111111111111111000000",
"10110100001111100001011100000010",
"11110110000100100011111011110011",
"10010001000100011000100000010000",
"00111110000100000001000100001010",
"01111111001111101111001110100111",
"00000100010000100010101111111111",
"00000100010000001001100100000000",
"01011001001111100000111000000000",
"00010001100010100001000111111111",
"00001001100100011001000010001010",
"11111111110000000000110100110110",
"00010110000000100000001011111111",
"00010001000010101001000100010001",
"00011000100010011000100000010000",
"00001001100100001001000101010110",
"10010001000000000000111101000000",
"11110110110011100011111010010000",
"00111110111111110100110100111110",
"00010000000100011111111100110000",
"10111000101011011001100010001001",
"11111111111010111100001010011111",
"00001001000010010000100110001001",
"11100100100011011000100000010000",
"10000010000000101111111111111111",
"00011110000010000100000001000110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"10010000000110010010001000000100",
"00001111000011110000111110010001",
"00001000000001010001100100011001",
"00101101110001101000010000010110",
"10010110101011001001011100000000",
"01000001010001100000010000001110",
"00001010001010100010110100000000",
"01000110000000000000011001000010",
"00000011010000000000000000110000",
"00000000001101110100011000000000",
"00010111000100010001101000010111",
"00010000000011100001111100101010",
"00111111010000100001110000110110",
"00001110000110010000100000000000",
"00000000010000010100011000000100",
"01000010000010100010101000101101",
"00110000010001100000000000000110",
"00000000000000110100000000000000",
"00010111000000000011011101000110",
"00010111000100010000111000011000",
"00000000000001010100001000101001",
"00000010010000001101011000001000",
"01001100110101110000101000000000",
"01000010000010100010101000101101",
"00110000010001100000000000000110",
"00000000000000110100000000000000",
"00010110000000000011011101000110",
"10001000000100000000001100001111",
"11111111101110100100000010011001",
"00001000010000100000101010001001",
"00000000001100010100011000000000",
"11111110000111010011111001010110",
"01000000010001100011110100011000",
"00000001000000000100011000001000",
"00001010101010000100011000010110",
"10101000010001100011110100000001",
"00001110000110010000001000001010",
"00000001000010101010100001000110",
"00000000000000100011110100000011",
"01000010001010100010001100111100",
"00101101010001100000000000000110",
"11111111111001100011111000000000",
"01001000000000000000010000111101",
"00001101010001000100110001001111",
"00000010111111111111111111100100",
"11101110101000100011111000000010",
"00001010100100010000100010010000",
"01001100100010010001000000010001",
"00000111010000100010101000101101",
"00110000010001100000100000000000",
"00000000000001000100000000000000",
"00000000010000010100011000010111",
"11111111101110100011111000010110",
"01010011000000000000010000111101",
"00111110010011100100011101001001",
"00001111000011111111111111010001",
"11110110010000100010110000100010",
"00000000000000010011110111111111",
"10101000010001100000100100100011",
"01000000010001100000001000001010",
"00000001000000000100011000001000",
"00111101000101110000111100010110",
"01010011001000110000000000000010",
"00111110000010011001000110010000",
"11010110001111101111111110000000",
"10010101001111100001000111111111",
"11111111110111010011111011111111",
"00010111100010010001000000001010",
"10010000100100010101011000100001",
"00000000000001110100000000001001",
"00111110000000000010000001000110",
"10101101100110001111111101110000",
"11110011110000101001111110111000",
"00000010001111011000100111111111",
"10010000001111100010001100000000",
"00010000010101100000100110010001",
"01111110001111101000100100010001",
"11110010001111100011110100000000",
"11101100001010000011111011111111",
"01010101000000000000010000111101",
"01010110010100100010111000101110",
"00111101111111111110111100111110",
"00101110010101010000000000000011",
"00001000100100011001000001010010",
"00101001000100000001011100001110",
"00100001000000000000000101000010",
"00111110100010010001000000010001",
"00001110010101101111111110011110",
"00111101111111111000011000111110",
"00101110010101010000000000000010",
"00111110111111111110001000111110",
"00000011001111011110101111110110",
"01010010001011100010111000000000",
"11111111111100000011111001010110",
"00101110000000000000001000111101",
"00100101001111100101011001010010",
"00000000000000010011110100000000",
"10010001000010001001000000101110",
"00001001010000100010101000001111",
"00001000100100000010000100000000",
"00001010001001100000111101010110",
"00010000000100011000100000010000",
"11111111011000000011111010001001",
"01001000001111100000111001010110",
"00000000000000100011110111111111",
"11011100001111100010111001000100",
"11101011101110000011111011111111",
"01000100000000000000010000111101",
"01010110010100100010111000101110",
"01010110111111110100010100111110",
"11111111001011010011111000001110",
"01000100000000000000001100111101",
"00111110010000110101001000101110",
"00001110010001001110101011011001",
"00000001111111111101100001000110",
"01010101000000000000010100111101",
"01010010001011100010111001000100",
"11111111111011000100011001000011",
"00000000000100100100011000000010",
"00000000000100100100011000011100",
"10111011010000100010110000010111",
"11111111111000000100011000000001",
"00000000010001100000111000000010",
"00001110001010100001011100000001",
"00001010010111001100011000011000",
"00010000000101100000001000010000",
"01001100010001100000000110001000",
"00011100001011000000010000001010",
"00001010010011000100011001010110",
"00000001010100110100001000000011",
"00000001000000001100011000001110",
"00000000111111110100011000000000",
"01000010000010100010110000101101",
"01010111000010000000000000001000",
"01000000110110110000110101000000",
"01000110000000000000000100111100",
"00101100001011010000000011111110",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"00101001010000000001000000000001",
"11111101010001100000000000000001",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000001000101100100000000010000",
"00000000111111000100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000010000001101000000",
"00101101000000001111101101000110",
"00001111010000100000101000101100",
"01000110000011100000100000000000",
"00001101000000011111111111011000",
"00000100000000000000111011110110",
"00000000111010100100000010111101",
"00000000111110100100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000001101011101000000",
"00101101000000001111100101000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000011000100",
"00101100001011010000000011111000",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"10110001010000000001000000000001",
"11110111010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000000100111100100000000010000",
"00000000111101100100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000010000101001001000",
"00000000000000001000101101000000",
"00101101000000001111010101000110",
"00001001010000100000101000101100",
"01001000010001100000100000000000",
"01000000000100000000000100001010",
"01000110000000000000000001111000",
"00101100001011010000000011110100",
"00000000000010010100001000001010",
"00001010010010000100011000001000",
"01100101010000000001000000000001",
"11110011010001100000000000000000",
"00001010001011000010110100000000",
"00001000000000000000100101000010",
"00000001000010100100100001000110",
"00000000010100100100000000010000",
"00000000000110110100011000000000",
"01000010000010100010110000101101",
"01000110000010000000000000001001",
"00010000000000110000101001001100",
"00000000000000000011111101000000",
"00101101000000000001101001000110",
"00001110010000100000101000101100",
"01001101010001100000100000000000",
"01000110010101100000001100001010",
"00010000000000110000101001001110",
"00000000000000000010011101000000",
"00101101000000000001100101000110",
"00001110010000100000101000101100",
"01001101010001100000100000000000",
"01000110010101100000001100001010",
"00010000000000110000101001001110",
"00001000000000000000111101000000",
"00000000000100000100011000001110",
"00000101010000100010101000010111",
"00001010010011100100011000000000",
"00001110100010000001000000000011",
"00010111000000010000000001000110",
"00000000001110000100001000101010",
"00000100000010100100111001000110",
"00011010000110100001101000011010",
"00010110000010010100000001000110",
"10001110000000100001110110010000",
"10011101100011101001110110011101",
"01011100001011010000001000010000",
"00001110000000000001101001000010",
"00000001100010000001000000011000",
"00101101000101100000001000010000",
"00000011010000100001111101011100",
"00001110001000010001011100000000",
"00010110000000100001000100001010",
"00001110000011101000111000000011",
"00001001100010001000100100001110",
"11111110001101010100000000001000",
"11011000010001100000111001000100",
"11000110001111010000000111111111",
"01010111100000101111111111010100",
"00000001111111111110010001000110",
"11001110000010011001000110010000",
"00010000110001101010110010010111",
"00000000110101101001110000000000",
"00001010001011000010110101010100",
"00001000000000000000010101000010",
"00000000000011100100000010011110",
"00101100001011010101010100000000",
"00000000000001010100001000001010",
"00000001010000001001100000001000",
"11010010101000100000100000000000",
"00101100001011010101001000000000",
"00000000000001100100001000001010",
"01000000100101111000111000001000",
"01010011000000000000000000001110",
"01000010000010100010110000101101",
"10011010000010000000000000000101",
"00001000000000000000000101000000",
"11111111111001001100011010100010",
"00010000000000100101101010000001",
"00011010100010000001000000010110",
"01000110111011000001100000111110",
"11000110000000011111111111101000",
"00111101100000011111111111010100",
"10000010111111111110010011000110",
"00000000000111000100101000010000",
"00001010001011000010110101010110",
"00001000000000000000010101000010",
"00000000000011110100000001010010",
"00101100001011010100111000000000",
"00000000000001010100001000001010",
"00000010010000000101001100001000",
"00010000010101000000100000000000",
"01010100000000000001110001010011",
"01000010000010100010110000101101",
"01010100000010000000000000000101",
"00000000000000000000111101000000",
"00001010001011000010110101010101",
"00001000000000000000010101000010",
"00000000000000100100000001010101",
"11000110010011110101011000001000",
"11000010100111000000000000010000",
"01011010000110000000000000000001",
"11111111111010001100011000000010",
"00010000000101100001000010000010",
"10110110001111100001101010001000",
"00000000000001100011110111101011",
"01010011010101000100010101010011",
"00111110010011110100111101001001",
"10010000000010010000100101010001",
"00000100000100001001100000000100",
"10011000000001000001000010011000",
"00010000100110000000010000010000",
"00100010001000000100111000000100",
"01000110000001000001000010011000",
"00100010001000000000000000010000",
"00000100100010000001000010011000",
"00100000000000000001100001000110",
"11111111000011110011111000100010",
"01000111000000000000011000111101",
"01001001010100110101010001000101",
"00011110001111100101010101001111",
"00000000000100000100011000000110",
"01000110111010000100001100111110",
"01000110000000100000100101001100",
"00010111000011110000010000000000",
"11101000011111110011111000001110",
"01111010001111100010001101001110",
"01110110001111100101011011101000",
"00000000000110100100011011101000",
"01010111111010000010011100111110",
"00111101000001011111100000111110",
"00000101111100110011111001010101",
"00000010000010010100110001000110",
"00000000001100000100001000101100",
"00111110000000000001000001000110",
"00000000010001101110100000010000",
"01010010001111100000111000000100",
"00111110001000110100111011101000",
"00111110010101111110100001001101",
"00011010010001101110100001001001",
"11100111111110100011111000000000"
)
,(
"00000010111111111101010001000110",
"11111111110101000100011001010101",
"00001001010011000100011000000001",
"11111111111110010100001000000010",
"00000001111111111101010001000110",
"00000010111111111101010001000110",
"00000010000010010100000001000110",
"00000010000010010100100001000110",
"01001100010001100000010000010110",
"00010111010101010000001000001001",
"01001100010001100010010101010110",
"01001000010001100000000100001001",
"01000110000110000000001000001001",
"01000110000111000000001111111111",
"10010001000000010000100101001000",
"01000110100010000001000000001010",
"01010111000000011111111111010100",
"00111101000001011000100000111110",
"01000101010010110000000000000100",
"00111110010101010011111101011001",
"00101101000011100000010101111101",
"00000000000001110100001000101100",
"11111111011111000011111000001000",
"10001101111111111111010001000000",
"00000010111111111111111111111100",
"11011010100101101101001110000010",
"00101101100111101000111010011100",
"00000000000010010100001000110110",
"00111110100110000000001100010000",
"11110010010000001111111101100010",
"10010111100011110000100111111111",
"10000101100011111001100110011001",
"00111110010101111000100000010000",
"00000011001111010000010101001001",
"01011001010001010100101100000000",
"00011110111111111011111100111110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"00000100001111010010001000000100",
"01010010010011110101011100000000",
"11010100110001100000100001000100",
"01001000010001101000001011111111",
"01001100010001100000000100001001",
"11010100110001100000000100001001",
"00000101001111011000000111111111",
"01010010010000010101000000000000",
"11010100110001100100010101010011",
"01001100010001101000001011111111",
"01001000010001100000001000001001",
"11000110010101010000001000001001",
"00111101100000011111111111010100",
"01000101010100100000000000001101",
"01010010010011110101010001010011",
"01001110010010010010110101000101",
"01010110010101000101010101010000",
"11000000001111100101010100001110",
"00000000000010100011110111111111",
"01000101010101100100000101010011",
"01010000010011100100100100101101",
"11101010001111100101010001010101",
"11111110101110010011111011111111",
"01010001000000000000010100111101",
"01011001010100100100010101010101",
"00000100110011110011111001010100",
"00111110110101100000100010010000",
"10010000000011101111111011010010",
"00001111111001110111101100111110",
"10010111110011101000111000000011",
"00000000000011111100001010101100",
"10011111101010011001100110001000",
"00011001000000000000010011000010",
"10011000000000000000000101000000",
"00011000000000000000110101000000",
"11000010101011001001011111001100",
"10001110100010100000000000000101",
"10011000000000000000000101000000",
"11000010100111111011100010101101",
"00010001000010001111111111001101",
"10010010001111100101100010001001",
"00000000000001100011110100000100",
"01001001010001100100010101010010",
"00111110010101010100110001001100",
"10101111001111100000010010000101",
"11111111111100000000110111111111",
"01010111000000010000001011111111",
"00111101000001000111100000111110",
"01000011010000010000000000000110",
"01010100010100000100010101000011",
"00001110100100000000100010010000",
"00001110000111010001011000000010",
"00101101000111010001011000000010",
"00000000010000110100001000111000",
"00001110000000101001110110010000",
"00000000000011100100001000011000",
"00010000000100010001011000010001",
"00000010100010000001000000011101",
"01000000000000000011101100111110",
"00010000000010000000000000101010",
"10011110111001000011011000111110",
"11001110100001001001100110001110",
"10011001100110011000111110100000",
"11010011100101101010001010000100",
"01000010100111001101101010010110",
"00010001000011100000000000001001",
"10010001000100011000100000010000",
"00001000000000000100110000111110",
"00000010100010000001000000010000",
"00010110000110100001101000011000",
"00001001111111111011100001000000",
"00000000000001100011110110001001",
"01000101010100000101100001000101",
"10010001010101100101010001000011",
"00100100010000000000100110010000",
"00000010100111011001000000000000",
"10010000100100010001011010010001",
"00100011010011100001000100000011",
"00010001000000110001000010011000",
"00100011000000000001000001000110",
"00010001000000110001000010011000",
"00100011000000000001100001000110",
"00010001000000110001000010011000",
"10001001000100010001000010001001",
"10011111101110001010110110011000",
"10001001111111111101011011000010",
"10010000001111010000101000001010",
"00010000100000101001000000001000",
"00000000100110100100001010011001",
"00001110000000100000111000011101",
"00001101000011110011011000011000",
"01111111111111111111111111111111",
"00101010000101110001000100011100",
"10000001010000100001110000011111",
"00001111000010101001000100000000",
"01010101000110101001000000010110",
"10000100100100000001100100100011",
"10011100000000001000000011000110",
"00001000100100001000101000010001",
"00000000001100001100001010101010",
"00011101000010110101001101001001",
"00000000111111110100011000000010",
"00101101010100110000000000011100",
"00001000010000100000101000101100",
"01000110000010000000100000000000",
"00001111010000000000000000111111",
"00101101010100100000000000000000",
"00000101010000100000101000101100",
"01000000100111100000100000000000",
"10011000000010000000000000000010",
"00000000100000000100011000010000",
"00000011000011110010001000011100",
"00011101000010110101010000011000",
"01000010010000111001101100011101",
"10010000000000100000000000000001",
"00010000000100010000100110010001",
"00100011010011100001000100000011",
"00010001000000110001000010011000",
"00100011000000000001000001000110",
"00010001000000110001000010011000",
"00100011000000000001100001000110",
"10001010000000110001000010011000",
"01000010000111000101010100010001",
"00011010000100010000000000000101",
"10001001000000110001100000010000",
"00010000000000010001000001010111",
"01000000000010000000111010001000",
"00001001000010001111111101100001",
"00000010000011100011110110001001",
"00001001100100001001000101010110",
"00011101000000000001101001000000",
"00001101000110000000001010010000",
"01111111111111111111111111111111",
"00011111001110000010110100011100",
"00000100010000100000111000001010",
"10001001100010000000101000000000",
"10001000000100000000100000111101",
"10011111101110001010110110011000",
"10001001111111111110000011000010",
"10010001001111010101011000001001",
"00001110100100000000100110010000",
"00001110000111010001011000000010",
"00101101000111010001011000000010",
"00000000100000100100001000111000",
"10010111110101111000001010010000",
"01110000110000100001110110101100",
"00001110000111100000111000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"00010110010100110001011000100010",
"10001000000100000001110001011010",
"00001111000010101001000100010001",
"01000010111111111001111100111110",
"00011110000011110000000001010010",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"01100011001111100010001000000100",
"00101011010111110000110111100101",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11100101010100000011111000100010",
"00010001111001011011101000111110",
"00000000001000110100001000101010",
"11100100110011100011111001000111",
"00111110000000000001100001000110",
"00111110000100001110010100010001",
"10010001100100000000011001001100",
"00000010000011110000111110010111",
"00010000000110100001101000011000",
"00010100001111100001011010001000",
"00000000000110100100011011100101",
"00010000111001001010111100111110",
"00001000100100001001100010001000",
"00011000000000100000111000001010",
"01000000000101100001101000011010",
"10001000000010011111111101111001",
"00001010001111011000100100010000",
"01101110011101010010000000000000",
"01101001011001100110010101100100",
"01010101011001000110010101101110",
"00000001111111111101010001000110",
"11111111110011000000110110111101",
"00001110000000100000001011111111",
"00000010000010100111110001000110",
"00001010100100010001011000011001",
"00001110000011101000100000010000",
"00011101000101100001110100000010",
"00001111000011110000100010010000",
"00111110000101110000111100010000",
"00001111000100001111110111001110",
"00101110001111100101011000010111",
"01011000010000100010101111111111",
"10001000000100000000100000000000",
"10000010111111111101010011000110",
"11000110111111111100010000111110",
"00000111100000011111111111010100",
"00000000001001100100001000101100",
"11111111111111111100110000001101",
"01000110000011100000001000000010",
"00011001000000100000101001111100",
"00010000000010101001000100010110",
"01010101000011110000111110001000",
"10010111001111100001101000011010",
"00011010000110100101010111111101",
"00000010000010101000000001000110",
"01000000111111101111010000111110",
"00000100001111100000000000011100",
"00101011111101110000110111100101",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11100100100001000011111000100010",
"00111110111001001110111000111110",
"00000001010000001110001100000100",
"01001111001111011000100000000000",
"00101010001010100010101000000000",
"00101010001010100010101000101010",
"01100001011001000010000000101010",
"01110011001000000110000101110100",
"01101011011000110110000101110100",
"01110010011011110110001100100000",
"01110100011100000111010101110010",
"01110100001000000110010001100101",
"01110101011011110111001001101000",
"01101001001000000110100001100111",
"01101001011101000110100101101110",
"01100011001000000110110001100001",
"00101100011001010110010001101111",
"01110010011011110110011000100000",
"00100000011100110110010101100011",
"01100101011100100010000001100001",
"01110010011000010111010001110011",
"00100000001000010010000001110100",
"00101010001010100010101000101010",
"00101010001010100010101000101010",
"11111111111111111100110000001101",
"10000100010001100000001000000010",
"01000110001011000000001000001010",
"00101100000000100000101010000000",
"00000000000011110100001000100010",
"11111111111111111111110000001101",
"01110100010001100000001000000010",
"01000110000011100000000100001010",
"01010110000000010000101010000100",
"00000001000010100101110001000110",
"00001010010011110100011001010111",
"11110000010001100101011100000011",
"00000100000011100011111000000000",
"00000010000010100101110001000110",
"01111100010001100000111100100010",
"01000110000011100000000100001010",
"00001010000000010000101001111000",
"00000000010010110100001000101100",
"11111111111111111100110000001101",
"01010001100100000000001000000010",
"01001111001111100001110100010000",
"11111110110100010011111011100000",
"00010001000111111001000000111000",
"00000010000010100111110001000110",
"00011100000001000001011000011001",
"00010001000000000000111101000010",
"00010110000000101000100100001110",
"11111111110011000000110100011101",
"01000000000000010000001011111111",
"01111000110001100000000000011101",
"01110100010001101000000100001010",
"11111100000011010000001000001010",
"00000001000000101111111111111111",
"10000100010001100101011010001000",
"00011101000000100000111000001010",
"00111110111000001110101000111110",
"01000111000000011110000100111110",
"01000110111000110001101100111110",
"01011110001111100000000000010100",
"00001010010111000100011011100011",
"00000100100101100011111000000010",
"00000010000010100111100001000110",
"00000000000110100100011000110110",
"11100011000000100011111000010110",
"00001010010011110100011001010110",
"00111110010101110011110100000011",
"00101100100100000000001111001101",
"10010001000000000110000101000010",
"00101101100010000001000000010110",
"00000000010110000100001000111000",
"00001110000111011000001010010000",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00010110001000100000010000011001",
"00011100010110100001011001010011",
"11100000100110010011111000001111",
"10010001000000000000101101000010",
"01010010100010010001000000010001",
"01000000111111001100000000111110",
"10001000000010000000000000101000",
"00001110000111100000111110011000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11100011001010000011111000100010",
"00000000001011011010001100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110111000110001010100111110",
"00001110000010101110001101111111",
"00011010000110100001100000000010",
"11111111101000110100000000010110",
"10000100010001100101011000001001",
"00010011110000101011010100001010",
"00001010011101000100011000000000",
"11111111111111000000110100000010",
"00001110000000010000001011111111",
"01000000001111100001110100000010",
"11100000100101000011111011100000",
"01110001001111100100011100000001",
"00000000000101000100011011100010",
"00010000111000101011010000111110",
"11101101001111100000111010001000",
"00011010010001100011011000000011",
"01000110010101010001011000000000",
"00111110000000011111111111010100",
"00001011001111011110001001011000",
"01101110011101010010000000000000",
"01101111011100110110010101110010",
"01100100011001010111011001101100",
"00100010010101010011110101001110",
"01000100000000000000001100111101",
"00111101010100100101001001001001",
"01001001010000100000000000000011",
"00000011001111010101010001001110",
"01001111001011110101011100000000",
"00000000000000110011110101010000",
"11000110010011110010111101010010",
"01000110100000101111111111010100",
"00001111000011110000101010011100",
"00001111100100000001011000000010",
"11000110101011000000100100000001",
"10011100100000100000101010100100",
"00111110000000000000001111000010",
"11010100110001100000000000001010",
"00000011001111011000000111111111",
"01010111001011110101001000000000",
"00000010000010100101100001000110",
"00000000000010100100001000110101",
"00001010101001000100011001010110",
"00111110010101110000111000000001",
"00111101000010001110000000010010",
"01001111010011000000000000000111",
"00101111010010010100101101000011",
"11111111110101000100011001001111",
"01000110000011100101011000000010",
"01000110000000110000101001001101",
"01000110000000010000101001011100",
"01000110000000011111111111010100",
"00110110000001000000101001001101",
"01000110111111111111100001000010",
"01000110000000101111111111010100",
"01000110000001000000101001001101",
"00100001000101110000000000011010",
"00000010000010100101110001000110",
"01000110000011100101011000010110",
"01000110000000110000101001001101",
"00001111000000010000101001011100",
"00000001111111111101010001000110",
"01010101010010000011110100001010",
"01000110000010011001000010010001",
"01010101000000100000101001010000",
"00001111000011110010000000010000",
"00001000010000100010110000011100",
"01010000010001100010001000000000",
"10001001000100000000000100001010",
"10101101100110000000100100111101",
"11100010110000101001111110111000",
"00111101010101111000100111111111",
"11111111010101110011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"01110101001111100100011100000001",
"10111010001111100100011111100001",
"10110110001111101001000011100001",
"00000000000110100100011011100001",
"00111110111000010110011100111110",
"01000010001010111111111101111011",
"10011011100110110000000000010011",
"00010000010101011001101110011011",
"00100010010101010001111100100000",
"00010000000010100101000011000110",
"00000001000100000001110000000010",
"11010100110001101000100010001000",
"00111110010101111000000111111111",
"01010101001111011111111100011001",
"11000110111111110001010000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"10000101001111100000100010010000",
"00011010000110100001101011111111",
"00011111001010010010001000011010",
"10010000000000000001110101000010",
"11100001001000100011111001000111",
"11100001011001110011111000010001",
"00111110111000010110010000111110",
"00011010010001101110000101110111",
"11100001000100100011111000000000",
"00100100001111101000100100010000",
"00000000000001000100000011111111",
"00001110000010100000101010001000",
"10000001111111111101010011000110",
"11111110110100110011111001010111",
"01000011000000000000101000111101",
"01000101010100110100111101001100",
"01001100010010010100011000101101",
"11111110101011100011111001000101",
"10100110001111100101010100100010",
"00111110010101100011110111111111",
"00001011001111011111111110100001",
"01000101010100100100001100000000",
"00101101010001010101010001000001",
"01000101010011000100100101000110",
"11111110101001110011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"11000101001111100100011100000001",
"00001010001111100100100011100000",
"11100001000111010011111011100001",
"00111110000000000001101001000110",
"11001100001111101110000010111000",
"11111111110101001100011011111110",
"10000010001111100101011110000001",
"00000000000010010011110111111110",
"01001110010001010101000001001111",
"01001100010010010100011000101101",
"01110010001111100101010101000101",
"11111111110101001100011011111110",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010100001110000010010000",
"11010010001111101110000011010101",
"00000000000110100100011011100000",
"00001101111000001000001100111110",
"00000010111111111111111111111100",
"01011010000101100101001100000010",
"11110000010001100100111000011100",
"00000000110100100011111000000000",
"11111110100001010011111000001000",
"11111100000011010000100010010000",
"00000010000000101111111111111111",
"00011100010110100001011001010011",
"00010000000000100001110110010000",
"10001000000100000000001010001000",
"10000001111111111101010011000110",
"11111110001001110011111001010111",
"01000100000000000000101100111101",
"01010100010001010100110001000101",
"01001001010001100010110101000101",
"00111110010101010100010101001100",
"11010100110001101111111000010101",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01001110111000000011001100111110",
"00111110111000000111100000111110",
"00011010010001101110000001110101",
"11100000001001100011111000000000",
"11111111111111111111110000001101",
"00010110010100110000001000000010",
"01000110010011100001110001011010",
"01110101001111100000000011110000",
"00101000001111100000100000000000",
"00001101000010001001000011111110",
"00000010111111111111111111111100",
"01011010000101100101001100000010",
"00000010000111011001000000011100",
"00010000000000101000100000010000",
"11111111110101001100011010001000"
)
,(
"11001010001111100101011110000001",
"00000000000011010011110111111101",
"01000101010011000100100101000110",
"01010011010011110101000000101101",
"01001111010010010101010001001001",
"00001001001111010000100001001110",
"01001100010010010100011000000000",
"01001001010100110010110101000101",
"00111110010101010100010101011010",
"11010100110001101111110110101001",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01001100110111111100011100111110",
"00111110111000000000110000111110",
"00011010010001101110000000011111",
"11011111101110100011111000000000",
"11000110111111011100111000111110",
"01010111100000011111111111010100",
"00111101111111011000010000111110",
"01001110010010010000000000001100",
"01000100010101010100110001000011",
"01001001010001100010110101000101",
"10010000100100010100010101001100",
"00011100000000001111000001000110",
"00010110000010010100000001000110",
"00010000000000010001110110010000",
"01010110100111011001110100000001",
"00010000100111010000111100010000",
"10001000000100000000000100000001",
"00000000000010000011110110001001",
"01001100010000110100111001001001",
"01000100010001010100010001010101",
"00011010000110100001110001000111",
"00010110000010010100000001000110",
"00111110010101010011110100000010",
"11010100110001101111110101000001",
"01000110010101011000001011111111",
"10010001000000011111111111010100",
"11111111101111100011111010010000",
"00111110010001110000100010010000",
"00111110010101001101111101011000",
"10001010000100011101111110011101",
"00010001110111111001100000111110",
"00000000110100100011111010001010",
"00111110000000000001101001000110",
"01011000001111101101111101000100",
"00010001000010001001000011111101",
"11000110100010010001000000000010",
"01010111100000011111111111010100",
"00111101111111010000100000111110",
"01001100010000100000000000000101",
"01010101010010110100001101001111",
"11000110111111001111110000111110",
"10010000100000101111111111010100",
"11111111111111000000110100001000",
"01010011000000100000001011111111",
"00010000000111000101101000010110",
"00111110000000001111000001000110",
"00001000100100001111111101110000",
"11011111000010100011111001000111",
"00111110000000000001011001000110",
"11110000010001101101111101001101",
"11011111010001110011111000000000",
"10000001001111101000101000010001",
"11010100010001100101010100000000",
"00011010010001100000000111111111",
"11011110111011100011111000000000",
"10010000111111010000001000111110",
"11111111111111000000110100001000",
"01010011000000100000001011111111",
"00010001000111000101101000010110",
"11000110100010010001000000000010",
"01010111100000011111111111010100",
"00111101111111001010100000111110",
"01000101010100100000000000001001",
"01000110001011010100010001000001",
"01010101010001010100110001001001",
"11000110111111001001100000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11110000010001101001000010010001",
"01000000010001100001110000000000",
"00011101100100000001011000001001",
"10011101000000010001000000000001",
"00001111000100000101011010011101",
"00000001000000010001000010011101",
"00111110010001111000100000010000",
"00111110010100111101111010011100",
"00111110000100001101111011100001",
"00111110000100011101111011011101",
"00011010010001100000000000011000",
"11011110100010100011111000000000",
"11111100100111010011111010001001",
"00010000000000100000100010010000",
"11111111110101001100011010001000",
"01001110001111100101011110000001",
"00111110010101010011110111111100",
"00111110000011101111110001001001",
"00100011010011101101111010111001",
"11011110101100110011111000001110",
"00111110000011100010001101001110",
"00100011010011101101111010101101",
"01010111110111101010100000111110",
"00111101111111000011000000111110",
"01000101010100100000000000001001",
"01001100001011010100010001000001",
"00111110010001010100111001001001",
"11010001001111101111111111010100",
"00111110010101010011110111111111",
"11010100110001101111110000011001",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"01001111110111100011011100111110",
"00111110110111100111110000111110",
"11011110001111101101111001111001",
"00000000000110100100011011111111",
"00111110110111100010011100111110",
"11010100110001101111110000111011",
"00111110010101111000000111111111",
"01010101001111011111101111110001",
"11000110111110111110110000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011110000010100011111001000111",
"11011110010011110011111001001101",
"00111110110111100100110000111110",
"00011010010001101111111110110001",
"11011101111110100011111000000000",
"11000110111111000000111000111110",
"01010111100000011111111111010100",
"00111101111110111100010000111110",
"01000101010100100000000000001111",
"01001001010100110100111101010000",
"01001110010011110100100101010100",
"01001100010010010100011000101101",
"10101110001111100101010101000101",
"11111111110101001100011011111011",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00010010010001101101110111001100",
"11011110000011110011111000000000",
"00111110110111100010001000111110",
"00011010010001101111111101110001",
"11011101101110100011111000000000",
"11000110111110111100111000111110",
"01010111100000011111111111010100",
"00111101111110111000010000111110",
"01000101010100100000000000001011",
"01000101010110100100100101010011",
"01001100010010010100011000101101",
"01110010001111100101010101000101",
"11111111110101001100011011111011",
"11010100010001100101010110000010",
"00011011000110110000000111111111",
"10001101001111100001101100011011",
"11011101111010010011111011011101",
"00111110000000000001101001000110",
"11010100110001101101110110000100",
"01010111010101101000000111111111",
"00111101111110110101000000111110",
"01000101010100110000000000001100",
"01001001010001100010110101010100",
"01000001010001000100010101001100",
"00111110010101010100010101010100",
"11010100110001101111101100111101",
"01000110010101011000001011111111",
"00011011000000011111111111010100",
"00111110000110110001101100011011",
"10110100001111101101110101011000",
"10011010001111100100100111011101",
"10010110001111100100110011011101",
"00000000000110100100011011011101",
"11000110110111010100011100111110",
"01010110100000011111111111010100",
"11111011000100110011111001010111",
"01010111000000000000101000111101",
"01000101010101000100100101010010",
"01001100010010010100011000101101",
"00000010001111100101010101000101",
"11111111110101001100011011111011",
"11010100010001100101010110000010",
"00111110010001110000000111111111",
"00111110010010101101110100100000",
"01111000001111101101110101100101",
"00000000000110100100011011011101",
"00001101110111010001001100111110",
"00000010111111111111111111111100",
"01011010000101100101001100000010",
"11110000010001100101001000011100",
"11111101011000100011111000000000",
"11111011000101010011111000001000",
"11111100000011010000100010010000",
"00000010000000101111111111111111",
"00011100010110100001011001010011",
"11000110100010000001000000000010",
"01010111100000011111111111010100",
"00111101111110101011110000111110",
"01010010010101110000000000001010",
"00101101010001010101010001001001",
"01000101010011100100100101001100",
"11111010101010110011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"11001001001111100100011100000001",
"00000000000100110100011011011100",
"00111110110111010000110000111110",
"00011010010001101101110100011111",
"11011100101110100011111000000000",
"11111111111111111111110000001101",
"00010110010100110000001000000010",
"01000110010011100001110001011010",
"00001001001111100000000011110000",
"10111100001111100000100011111101",
"10001101000010001001000011111010",
"00000010111111111111111111111100",
"11011010100101101101001110000010",
"00000010000111010001000010011100",
"10001001000100010000001000010000",
"10000001111111111101010011000110",
"11111010010111110011111001010111",
"01000110000000000000101100111101",
"00101101010001010100110001001001",
"01010100010000010101010001010011",
"01010110000010000101001101010101",
"01000111000000000000110000111101",
"01000110001011010101010001000101",
"01000100010001010100110001001001",
"01010101010001010101010001000001",
"11000110111110100011110000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011100010110100011111001000111",
"11011100100111110011111001001001",
"00001110000010011001000010010001",
"00001110110111001001100000111110",
"10010010001111100010001101001110",
"11011100101001010011111011011100",
"00001110100010010001000000010001",
"00001110110111001000100000111110",
"10000010001111100010001101001110",
"11011100100101010011111011011100",
"00111110000000000001101001000110",
"01000100001111101101110000110000",
"11111111110101001100011011111010",
"11111010001111100101011110000001",
"00000000000010100011110111111001",
"01010011010101010100110001000110",
"01001001010001100010110101001000",
"00111110010101010100010101001100",
"11010100110001101111100111101001",
"01000110010101011000001011111111",
"01000111000000011111111111010100",
"00111110110111000000011100111110",
"00111110000011101101110001001101",
"01001110000011101101110001001001",
"11011100010000110011111000100011",
"10010001110111000101011000111110",
"00111110000000001111000001000110",
"00001000100100001111110001010000",
"00111110000000000001101001000110",
"11111100001111101101101111101000",
"10010001100010100001000111111001",
"00010000000000100001000100001010",
"11111111110101001100011010001001",
"10101010001111100101011110000001",
"00000000000010110011110111111001",
"01000001010011100100010101010010",
"01000110001011010100010101001101",
"01000110010001010100110001001001",
"10101001001111100000000000010000",
"00010001010001100011110111111111",
"11111111101000100011111000000000",
"01000001000000000000110100111101",
"01001100010011110101001101000010",
"00101101010001010101010001010101",
"01000101010011000100100101000110",
"11111001011110110011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"10011001001111100100011100000001",
"11011110001111100101001011011011",
"00000000000000000000110111011011",
"11011000000011010000001100000000",
"00000010000000101111111111111111",
"01000000000010011001000010010001",
"00000010000100000000000000100101",
"00011001000011100001111000001110",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"11010000001111100000101000011110",
"00001110000111010001000011011011",
"11011011110010010011111001010010",
"11000100001111100101001000011101",
"00011010000110100101001111011011",
"10101101100101100000100010010000",
"11010101110000101001111110111000",
"00011010010001101000100111111111",
"11011011010100100011111000000000",
"10000001111111111101010011000110",
"11111001000111110011111001010111",
"01000101000000000000110000111101",
"01001001010100100101010001001110",
"01000110001011010101001101000101",
"11000110010001010100110001001001",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011011001011100011111001000111",
"11011011011100110011111001001011",
"00111110000000000001101001000110",
"11010100110001101101101100100100",
"00001110001111011000000111111111",
"01000001010001010101001000000000",
"01000011010010010100010001000100",
"01001110010011110100100101010100",
"11000110010110010101001001000001",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011011000000100011111001000111",
"11011011010001110011111001010001",
"00111110110110110100010000111110",
"00011010010001101101101101000001",
"11011010111100100011111000000000",
"10000001111111111101010011000110",
"01010000000000000000010000111101",
"11000110010001010100011101000001",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011010110110100011111001000111",
"00111110000000000001011101000110",
"00011010001111101101101100011101",
"00000000000110100100011011011011",
"11000110110110101100101100111110",
"00111101100000011111111111010100",
"01010100010000010000000000000101",
"01010101010110010101100000101101",
"11000110111110001001000000111110",
"01010101100000101111111111010100",
"00000001111111111101010001000110",
"11011010101011100011111001000111",
"00111110000000000001110001000110",
"00011010010001101101101011110001",
"11011010101000100011111000000000",
"10000001111111111101010011000110",
"11111000011011110011111001010111",
"01000011000000000000110100111101",
"01000111010011100100000101001000",
"01000001010010000100001101000101",
"01010100010001010101001101010010",
"11111000010110110011111001010101",
"10000010111111111101010011000110",
"11111111110101000100011001010101",
"01111001001111100100011100000001",
"00000000000111010100011011011010",
"01000110110110101011110000111110",
"01101101001111100000000000011010",
"11111111110101001100011011011010",
"00111010001111100101011110000001",
"00000000000010100011110111111000",
"01000011010001000100010001000001",
"01001111010100110100111001001111",
"00111110000011110100010101001100",
"00100100010000100000100111000101",
"01000010001101010000111100000000",
"00000010000111010000000000001100",
"00010110000000000001000001000110",
"10001011001111100000111100000010",
"00001100010000100011011011010111",
"00011101000010001001000000000000",
"00000010000101100101011000000010",
"11100000010000001000100000010000",
"00000010010000000000100011111111",
"00111101010101100000100100000000",
"01010101010100110000000000001010",
"01001110010011110100001101000010",
"01000101010011000100111101010011",
"00001001100010110011111000001111",
"00001111000000000010000001000010",
"00000110010000100011010100001110",
"00111110000011110000100000000000",
"01000010001010110000000000100100",
"00001001100100010000000000001100",
"00010110010011100000001000011101",
"01000000100010000001000000000010",
"00001010000010101111111111100101",
"00001001000000000000001001000000",
"00000000000010100011110101010110",
"01010100010100110100111001001001",
"01000101010000110100111001000001",
"00001111000011110100011001001111",
"00101011111111111000101100111110",
"00001000000000000010010101000010",
"00001100010000100011010100001111",
"01000110000000100001110100000000",
"00000010000101100000000000010000",
"11010111000110000011111000001111",
"00000000000011000100001000110110",
"00000010000111010000100010010000",
"00010000000000100001011001010010",
"11111111111000000100000010001000",
"00000000000000100100000000001000",
"00000110001111010000101000001010",
"01010011010000010100001100000000",
"10010000010011110101010001010100",
"01000010001101011001000000001000",
"00000010100111010000000000010101",
"00100100000000100001000000001111",
"00001111001101100001110000010001",
"00000110010000100001110000110110",
"10011101100111010001100100000000",
"00001010111111111110110101000000",
"00000000000001000100001000001110",
"00000010000111010001000000001000",
"00001110100100010011110110001001",
"00111110010110101000100000010000",
"01000010001101011111111111010001",
"00001010000010100000000000000011",
"11101111000011010000100010111101",
"00011110000001000000000000110110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"11011011001111100010001000000100",
"11101101111010000011111011011001",
"00000000001101101110001100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00011101110110011100010100111110",
"00000000000100000100011000000010",
"00001110000111100000001000010110",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11011001101100000011111000100010",
"00000000001101101101011100001101",
"00011001000011100001111000000100",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110110110011001110100111110",
"00001010001111011101100000100000",
"01101111011011100010000000000000",
"01101111011001100010000001110100",
"00001010011001000110111001110101",
"01100110011011110010000000000000",
"01100001011011000110001100100000",
"00001100001000000111001101110011",
"01101110011011110110001100000000",
"01110101011100100111010001110011",
"01110010011011110111010001100011",
"01010011000000000000110100100000",
"01000011010100100100000101000101",
"01000101010011010010110101001000",
"01000100010011110100100001010100",
"00010001100100010000100010010000",
"00000000000111010100001010001010",
"00111110000011100000100010010000",
"00110101000111000000100001010001",
"01010010000000100001110100001111",
"00001111000011110000001000010110",
"00000101010000100001110000110110",
"01000000000010100000101000000000",
"00010000000010011111111111101101",
"00110110001111100000111110001000",
"01011001010000100001111100001000",
"00111000010111010000110100000000",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11011001001001000011111000100010",
"00001101111011010011000100111110",
"00000100000000000011100000111011",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"00111110000100001101100100001110",
"11100011000011011110110100011010",
"00011110000001000000000000110110",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"11110111001111100010001000000100",
"00000010000111010001000011011000",
"00010110000000000001000001000110",
"00011001000011100001111000000010",
"00001111001000000100111000000100",
"00100010000001000001100100011001",
"00111110110110001110000100111110",
"00111110000011111101011101100100",
"00110010010000100000011111010101",
"00110101110110100000111100000000",
"00001111000000000001111101000010",
"01001010000000100001110100001111",
"00111110000100000000001000010110",
"01000010001101011111111010100001",
"10010000100010010000000000000110",
"00111101000010100000101000001000",
"01010110000000100001110100001000",
"01000000100110110000001000010110",
"10010000000010001111111111011101",
"01001110000000100001110100001000",
"10001001000100000000001000010110",
"00001101111111111100011101000000",
"00000100000000000011100001011101",
"00000100000110010000111000011110",
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"10011111001111101101100010010010",
"00110110111000110000110111101100",
"00001110000111100000010000000000",
"00100000010011100000010000011001",
"00000100000110010001100100001111",
"11011000011111000011111000100010",
"01000110000000100001110100010000",
"00000010000101100000000000010000",
"00000100000110010000111000011110"
)
,(
"00011001000011110010000001001110",
"00111110001000100000010000011001",
"00100110000011011101100001100110",
"00011110000001000000000000111000",
"01001110000001000001100100001110",
"00011001000110010000111100100000",
"01010011001111100010001000000100",
"00111110100010000001000011011000",
"11010001001111101110110001011110",
"00000000000100110011110111010110",
"01110100011011110110111000100000",
"01110101011011110110011000100000",
"00100000001011000110010001101110",
"01100100011011100110000101101000",
"00100000001000000110010101101100",
"01100110011011110010000000000000",
"01100100011011100111010100100000",
"01101110011010010110011001100101",
"01101111001000000110010001100101",
"01100011011001010110101001100010",
"01110100011000010010000001110100",
"01100100011001000110000100100000",
"01110011011100110110010101110010",
"01101101000000000000011100100000",
"01101111011010000111010001100101",
"00000000000010110010000001100100",
"01000011010001010101100001000101",
"00101101010001010101010001010101",
"11000110010101110100010101001110",
"00110101100000101111111111010100",
"01000110000000000100010001000010",
"10010000000000100000101010010100",
"00001010100010000100011000011101",
"00010000010000100010101100000010",
"11101000010001100000100000000000",
"00000110011110110011111000000011",
"00000001000011110100110100001000",
"00001010100010000100011000001110",
"10000100001111101001000000000001",
"00001010001110000010110100001000",
"00010000000000000001000001000010",
"11101000010001100000111110001000",
"11000111001111100001011000000011",
"01000110100100000000100000000111",
"01000110000000010000101010001000",
"00010001000000010000101010010100",
"00000010000111011000100100010000",
"00001000000011100000000100010110",
"10000001111111111101010011000110",
"01000101000000000000111000111101",
"01010101010000110100010101011000",
"01001101001011010100010101010100",
"01001111010010000101010001000101",
"11111111110101001100011001000100",
"01000110000110100001101010000010",
"01010010000000100000101010010000",
"00000100010000100010101000101101",
"00010000000010101001000100000000",
"00010110100100000000100010001000",
"00000010000010101000110001000110",
"00000000000100000100001000101011",
"00000011111010000100011000001000",
"00001000000001100001000000111110",
"00001110000000010000111101001110",
"00000001000010101000110001000110",
"00001000000110010011111010010000",
"01000010000010100011100000101101",
"10001000000100000000000000010000",
"00000011111010000100011000001111",
"00000111010111000011111000010110",
"10001100010001101001000000001000",
"10010000010001100000000100001010",
"10001001000100010000000100001010",
"10000001111111111101010011000110",
"01010011000000000000100100111101",
"01001111010011000100110001000001",
"01000101010101000100000101000011",
"10000010111111111101010011000110",
"10000010000010101000110011000110",
"10010000010001101000001010011101",
"00101101000011110000001000001010",
"00000000000010010100001000111000",
"00010000000011110101011000011101",
"11110010010000000000000100010110",
"01000110000010011000100011111111",
"11000110000000010000101010010000",
"00111101100000011111111111010100",
"01000001010101100000000000001001",
"01000011010011110100110001001100",
"11000110010001010101010001000001",
"00001111100000101111111111010100",
"00001010100110000100011000110110",
"00001101010000100001110000000010",
"00000010000011100000111100000000",
"01000010001011000001011101010101",
"00001111010101000000000000000011",
"10001100010001100000100000000001",
"00000010000111010000001000001010",
"11010100110001100000000100010110",
"00000111001111011000000111111111",
"01010100010001010101001100000000",
"01010000010011110101010001010110",
"10000010111111111101010011000110",
"00001010011010000100011001010110",
"10011000010001100101011100000001",
"01000110010101010000000100001010",
"01010110000000011111111111010100",
"10010000000000101011101000111110",
"00010001000010011000001010010001",
"10010001010101101000100100010000",
"00000010000011100000100110010000",
"01001110000110100001101110010000",
"01001011010000100010110000010111",
"00100010010101000001000000000000",
"00001000100100000000000100001111",
"00000010000111010001000000011000",
"01001100001111100001000000010001",
"01010110000110110001101100000111",
"01000000000010011001000010010001",
"00010000000011110000000000101000",
"00000010000101100001101000011010",
"01000010000111000101010100001111",
"00001111001101010000000000000101",
"00110101000010100001110000000010",
"00010111010101010000001000001111",
"00001011010000100001110000101100",
"11111111110101001100011000000000",
"00000001000011110101010010000010",
"10000001111111111101010011000110",
"10111000101011011001100000001000",
"11111111110100101100001010011111",
"10001000000100000000100110001001",
"00010111010101001000100000010000",
"00000001000001010100001000101100",
"00010000000110000000100010010000",
"01010110000011100000001000011101",
"00001111001101010000001000010110",
"00101100000101110101010100000010",
"00000000000010110100001000011100",
"10000010111111111101010011000110",
"11000110000000010000111101010100",
"00001000100000011111111111010100",
"00000010000101100101001000001110",
"01010101000000100000111100110101",
"01000010000111000010110000010111",
"11010100110001100000000000001011",
"00001111010101001000001011111111",
"11111111110101001100011000000001",
"01001110000011100000100010000001",
"00001111001101010000001000010110",
"00101100000101110101010100000010",
"00000000000010110100001000011100",
"10000010111111111101010011000110",
"11000110000000010000111101010100",
"00001000100000011111111111010100",
"00000000000101001100011010010000",
"10001101100011101000001010010110",
"00000000000000001111111111111111",
"00000000011001011100001010011100",
"00000000001000000100011000001110",
"01000110000011110000001000010110",
"00000010000101100000000000101000",
"01010010000000100000111100110101",
"01000010000111000011011000010111",
"11010100110001100000000001001011",
"00001111010100101000001011111111",
"11111111110101001100011000000001",
"11111111000011010001000010000001",
"00011100000000000000000011111111",
"01000110000100000011100000011001",
"01010000001000110000000000010000",
"01000010001000100011100000010111",
"00000010000111010000000000101011",
"10010000100100010101011000001111",
"00000000000110100100000000001001",
"00001111001101010000001000001110",
"00101100000101110101010100000010",
"00000000000010110100001000011100",
"10000010111111111101010011000110",
"11000110000000010000111101010100",
"00001000100000011111111111010100",
"10111000101011011001100000011101",
"11111111111000001100001010011111",
"00101110010000000000100110001001",
"00000000000110000100011000000000",
"01010110000000100000111000010110",
"01000000000010011001000010010001",
"00001110000111010000000000011010",
"00000010000011110011010100000010",
"00011100001011000001011101010101",
"11000110000000000000101101000010",
"01010100100000101111111111010100",
"11010100110001100000000100001111",
"10011000000010001000000111111111",
"11000010100111111011100010101101",
"00001000100010011111111111100000",
"11010100110001101000100100010001",
"00001111010100101000001011111111",
"11111111110101001100011000000001",
"10011000000111010001110110000001",
"11000010100111111011100010101101",
"00001000100010011111111010010100",
"11111110011111110100001000101100",
"00001111000000010011101000111110",
"10010000100100010101011000000010",
"01010101000000100000111000001001",
"00000101010000100010110000010111",
"10110010001111100000111000000000",
"00011101000111010000100000000100",
"10011111101110001010110110011000",
"10001001111111111110101011000010",
"11111111110101000100011000001001",
"01000110010101100000100000000010",
"00111110000000010000101010011000",
"00000010000011110000000100001111",
"00001001100100001001000101010110",
"00001111010011100000001000001110",
"00000000000001110100001000011100",
"00000001000011110001110001011001",
"01010000000000000000100001000000",
"00000000000000110100001000011100",
"00011101000000010000111101010101",
"10111000101011011001100000011101",
"11111111111000001100001010011111",
"11010100110001100000100110001001",
"00000010001111011000000111111111",
"11000110001000010101011000000000",
"00111110100000101111111111010100",
"00111110100100000000000011110100",
"11111100000011010000011000101010",
"00000010000000101111111111111111",
"00010000001000000001000001010101",
"00011010000101110101001110001000",
"00111110000101100001101000011010",
"01100000010001100000011000101111",
"00010000000000011001000000001010",
"00111110000000010001110110001000",
"11010100110001100000000001001001",
"00001010001111011000000111111111",
"01010010010000010100110100000000",
"01010111010100110010011001001011",
"01010010010100000100010101000101",
"00001001111101010000010000111110",
"11111111101110110011111000000010",
"01000011000000000000100000111101",
"01010100010000010100010101010010",
"11000110010011010100110101000101",
"01000110100000101111111111010100",
"00110101000000100000101001100000",
"00001110000000000000011101000010",
"11111111111111111111110000001101",
"00010111000011100000000100000010",
"00001010011000000100011000001110",
"10001000000100000000000110010000",
"11010100110001100000000100011101",
"01000110001111011000000111111111",
"00011101100100000000101001100000",
"00000010100010000001000000000010",
"00000000001101010100001000110101",
"00011101000111010000111100001111",
"01010101000011101001000100000001",
"00001110000101100010000000010000",
"00010111010100111000100000010000",
"00000000010100010011111000011010",
"00001111000000010000111100001111",
"00001000000000010001110100001111",
"01010110000000010000111101010110",
"01001100000000010001110100001111",
"00000010001110000011111000001111",
"11111110010001100001110100011101",
"00000000001101010011111000000000",
"00001010011010000100011001010110",
"00001001001111010000100100000001",
"01001100010001010101001000000000",
"01000101010100110100000101000101",
"10010001010101100100110101001101",
"00001011010000000000100110010000",
"00001111000000100000111100000000",
"00001000100100000001110100000001",
"10011000100010000001000000011101",
"11000010100111111011100010101101",
"00001001100010011111111111101111",
"00001010011000000100011000111101",
"00011101000111010000111000000010",
"10010000100100010101011000111101",
"00000000000001010100000000001001",
"00011101000000010000111101010110",
"10011111101110001010110110011000",
"10001001111111111111010111000010",
"00100000110001100011110100001000",
"10001111100011111101011000000000",
"00010000010101011001101110010110",
"00001010010110110010110100100000",
"00010001000000000000111101000010",
"00010000000010001001000010001010",
"10010001100010100001000110001000",
"01000000100010000000100110010000",
"00010001100010100000000000000001",
"00111000000101110001100000010000",
"11111111110110100100001000011111",
"00010111001000000001000001010101",
"00010110000100000010000101011100",
"00101101010100010011110110001001",
"00000010010000100000101000101010",
"11000110001111010000100000000000",
"10011101000100000000101001100000",
"10000010000010001001000010000010",
"00010111000100010000111000011001",
"00011010000110100001101000100001",
"00100000000100010101010100010000",
"00001110100100010001011000010110",
"00010001000011100000001000011101",
"00100000000100000101010100010111",
"00010000010000100010110000100100",
"00000010000011100000100000000000",
"01010101000101110001000100001110",
"00101100001001000010000000010000",
"00001000000000000000001001000010",
"00011101100100000000111101010110",
"00000010100010000001000000000010",
"00110110000011110011011000010111",
"00000000001011000100001000011100",
"10001000000100000000111010010001",
"00001110000000101100000000111110",
"00010000010101010001011100010001",
"00010110000100010010010000100000",
"00001111001000000001000001010101",
"00001000000000000010000100111110",
"00010000010101010001011100010001",
"00010001000111000001111100100000",
"00011010010101000000111100010110",
"00011000000100000001011100011010",
"00001110000000100110011000111110",
"10001001100010000000100000001001",
"01001100000000000000010100111101",
"01000010010100110100110101000100",
"01100000110001101001000010010001",
"10000010100111010001000000001010",
"00001111100000100000100010010000",
"01000110000000000100001101000010",
"00001000000000101111111111010100",
"00101101010100110000001000001110",
"01000110000011110000101000111000",
"00101010000101110000000000100000",
"00011011010000100010110000011100",
"00011101000011100000100000000000",
"01010101000100000000001000011101",
"00001111000101100010000000010001",
"00011010001000010001011100010001",
"10010001000101100001101000011010",
"01010010001111101001000100001010",
"10001001000100010001000000000010",
"11111111110101000100011001010101",
"10010000110101011001000100000001",
"10010110000100001010000000001001",
"01000000100010000001000000010111",
"10001001000010011111111110111001",
"00001111100010010001000000010001",
"01000110000000000101111101000010",
"00001000000000101111111111010100",
"00101101010100110000001000001110",
"01000110000011110000101000111000",
"00101010000101110000000000100000",
"00000000001100110100001000011100",
"00011101000011111001000110010000",
"10000101001111100000111100000010",
"00010010010000100011010100000000",
"00111110000011110001000100000000",
"00110101000010100000000010101010",
"10010000000000000000100001000010",
"00011101000011110001110100011101",
"00001010100010000001000000000001",
"00000000000010100100001000110101",
"00010001010101010000111100010000",
"00111110001000000001011101010100",
"10001001000010001111111001110000",
"00001000000000000000010101000000",
"00000010000111010001110100001110",
"11111111110101000100011001010101",
"10010000110101011001000100000001",
"10010110000100001010000000001001",
"01000000100010000001000000010111",
"01000110000010011111111110011101",
"00001000000000101111111111010100",
"00001010011000001100011000111101",
"11010101000100001000111010000010",
"10010110101000001000001010001111",
"00001111001101100000001000001110",
"00011100001010100001011100010000",
"01010100000000000000011101000010",
"01000000000101100001101000011010",
"00010000000011101111111111101110",
"00010111010000100010110000010111",
"00000010000100010101010100000000",
"00111110000011110010000010010000",
"01010101000011101111111100010010",
"00100000000101110101010000010000",
"00010000111111100011101000111110",
"00000001000100010001100010001000",
"01100000110001100011110110001001",
"10000010100111010001000000001010",
"00010000100000100000100010010000",
"00010110001000000001000101010101",
"00100001000101110001000100001111",
"00011010000110100001101010010000",
"00001111001101100001000000010110",
"01000010000111000010110000000010",
"00011010010101000000000000001000",
"01000000100110010001011100011010",
"00000010000111011111111111101111",
"00111101100010011000100000001010",
"10000010100111011001110110010000",
"00010000000010100110000011000110",
"00001000100100001000001010011101",
"00010001010101010000111110000010",
"00010001000101100001000000100000",
"00011010000101110001000110001010",
"10010001000101100001101000011010",
"00111110000011110000111100001010",
"10001010000100010000000101000001",
"10010000100100011000101000010001",
"00010001100010000001000000001001",
"01000010001101100001011110010001",
"00011010010101000000000000010110",
"00001111100110010001011000011010",
"00010000010101010001011100010001",
"00010110000100010010010000100000",
"11101000001111100001000000001111",
"11111111111000010100000000000000",
"00010000000000011001000000001000",
"10010000001111011000100110001001",
"01111101001111100000111000001000",
"00001000010000100010101111111111",
"11001111001111100000100000000000",
"01110001001111100000111011111010",
"00001001010000100010101111111111",
"00111110000011100000100000000000",
"00111110000011101111110111100100",
"01000010001101011111111101100100",
"10001011001111100000000000001100",
"01000010001101010000111011111111",
"00001111000100000000000000000100",
"00001010100010000000000100011101",
"00000000000110110011111000111101",
"00000000000001110100001000101011",
"00000000000100000100011000001111",
"00111101000010000000000100001111",
"01000101010000100000000000001101",
"01010010010001100101010001010011",
"01001100010000100100010101000101",
"00110101010010110100001101001111",
"11000110000000000101000001000010",
"01001011100000101111111111010100",
"00001110000111000101101000010110",
"00000010000010100110100001000110",
"00001010011010000100011000010110",
"11111101011000100011111000000001",
"00110101111111101101101000111110",
"00001111000000000001001101000010",
"11111111100010110011111000001111",
"00000000000010010100001000110101",
"00011101000011110001110100011101",
"00000001000011110101010100000001",
"00001010100100010000101000001110",
"00001111001101101000100000010000",
"00010010010000100001110000110110",
"00000010000111010000111000000000",
"00011010010101000000111101010101",
"01010100000000100001011100011010",
"00010111010101000010000000010111",
"11000110111111010001011000111110",
"00101011100000011111111111010100",
"01000001000000000000100000111101",
"01000011010011110100110001001100",
"01010101010001010101010001000001",
"01000110111011100110000000111110",
"00010111000000100000101001100000",
"10101100100111001100111110010000",
"10010000000110110001101100011011",
"01010101000110011001110010111000",
"00000010000010100110010001000110",
"00010111001000000001011101010011",
"00011100100010000001000000101010",
"11101110001111110011111001010111",
"01001101000000000000011000111101",
"01001111010011000100110001000001",
"10010000000010001001000001000011",
"10000010100111011001000010000010",
"00000001000111010000111100001111",
"00000011010000100010110000010001",
"00000001000011110000111100000000",
"00011101000011110001000000001000",
"00000001000011110101011000000001",
"00000000000000110100001000010000",
"10001001000000010001000000001110",
"10011101100111010000100010010000",
"00000000000010110011110110000001",
"01000100010011100100000101001000",
"01000001010101100100010101001100",
"10010001010001000100100101001100",
"10000010100111011001000110000010",
"00000000000001100100001000010000",
"01000000000000010001000000010001",
"00001111000100010000000000000011",
"00000111010000100001000100000001",
"00011101000100010001000000000000",
"00000000000001000100000000000001",
"00000001000111010000111100010000",
"11000110001111010000100110001001",
"00001110100000101111111111010100",
"00001111111111110111000000111110",
"00011100001101100000001000011101"
)
,(
"00000000011010100100001000001110",
"00001111010101100000100010010000",
"00001010011000001100011000000001",
"10010000100000101001110100010000",
"00001110110101101000001000001000",
"01001110000000101001000000011101",
"01010101000100001000000100010111",
"00001111000101100010000000010001",
"00010111100100010001000100000010",
"00011010000110100001101000100001",
"00010111000100010000111100010110",
"00100100001000000001000001010101",
"00000010000011100001011000010001",
"00001010001110000010110101010011",
"00000000001000000100011000001111",
"00001010000111000010101000010111",
"00011101000111010000111100101100",
"00101100000101110001000000000010",
"00000000000110010100001000011100",
"11111111011111110011111000001111",
"01010101000101110001000100001111",
"00011100000111110010000000010000",
"00001010100100010001011000010001",
"01001110100010000001000000001010",
"11000100010000001001100000010111",
"10001000000100000000100011111111",
"10001001111111110010111000111110",
"11000110000010101000100000010000",
"00111101100000011111111111010100",
"11111110111100110011111000001111",
"11000110000000001001101101000010",
"01010011100000101111111111010100",
"00001111000111000101101000010110",
"00011010010101000000001000011101",
"01010101000000100001011100011010",
"00010111010011100010000000001111",
"00111000001011010000111100001010",
"10010001000000000000010001000010",
"00001000100010000001000000001010",
"01011010000000010000010100111110",
"01000010001110000010110100011100",
"00001010100100010000000000000100",
"00011011000010001000100000010000",
"00001111000010001001000000011011",
"11111100000011010000001000011101",
"00000010000000101111111111111111",
"01011010000101100101001110010000",
"00011010000110100001000100011100",
"00010100001111100001011001010011",
"00000000000000000000000000000001",
"11111011100000100011111000010001",
"01010101000011111000001010010001",
"00011110001111100000000100001111",
"00010110010011100000100011111111",
"00001111111110111010101100111110",
"11011010001111100000111100001111",
"00001001010000100011010111111101",
"00001111000111010001110100000000",
"00001111000100000000000100011101",
"10001000000010100000111000000001",
"10001000000100000000101010010001",
"00011100001101100000111100110110",
"00010000000000000000110001000010",
"00011100010110100001011001010011",
"00010001000000100001110100001111",
"10001101111110110100011100111110",
"00000010111111111111111111111100",
"11000110001011001000100010000001",
"01000000100000011111111111010100",
"00111110000010100000000000000100",
"00000100001111011111110111010011",
"01000101010100100100011000000000",
"11111111110101001100011001000101",
"01000010001111100000111010000010",
"00000000000101000100001011111110",
"00011010010101000000001000011101",
"01010101000000100001011100011010",
"10001000000100000000101010010001",
"00011010000110100101010000100000",
"00000000000000100100000000010111",
"11010100110001100001011100001110",
"00000110001111011000000111111111",
"01010011010001010101001000000000",
"11000110010001010101101001001001",
"00001110100000101111111111010100",
"01000010111111100001010000111110",
"00000010000011100000000000000101",
"00001000000000010000111100011000",
"10000001111111111101010011000110",
"01000001000000000000111000111101",
"01000011010011110100110001001100",
"01000100010001010101010001000001",
"01011010010010010101001100101101",
"11111111110101001100011001000101",
"11101110001111100000111010000010",
"00000000000100000100001011111101",
"00010111010101010000001000001110",
"00001111001001010101011010010000",
"00000011110000101010110000000001",
"11111110011000110011111000000000",
"11111111110101001100011000001000",
"00000000000011000011110110000001",
"01010010010000110100111001001001",
"01010010010001010100011001000101",
"01000101010000110100111001000101",
"11111111111111111101100000001101",
"11111100000011010000001000000010",
"00000010000000101111111111111111",
"00000000000011000011110100010111",
"01010010010000110100010101000100",
"01010010010001010100011001000101",
"01000101010000110100111001000101",
"11111111111111111111110000001101",
"00010110010100110000001000000010",
"11111100000011010001110001011010",
"00000001000000101111111111111111",
"01010101000000000000011000111101",
"01000101010100110101010101001110",
"11111111111111000000110101000100",
"00010110000000100000001011111111",
"11111111111111111111110000001101",
"00000101001111010000000100000010",
"01001001010011000100000100000000",
"00111110010001110100111001000111",
"00010101010001101100111000001000",
"11001110010010110011111000000000",
"00111110111111111010100100111110",
"01000110010101011110111110000100",
"00011001000000100000101001100100",
"01111001001111100001101000100000",
"00000000000000000000110111101111",
"11001100000011010000010000000000",
"00000010000000101111111111111111",
"11101111011010100011111000010111",
"00111110000000000001101001000110",
"00000101001111011100110111011100",
"01001100010011000100000100000000",
"00111101010100000101010001001111",
"00010000001111010001110001010011",
"01001001010100100101010000000000",
"01010010010001010100011101000111",
"01010011010110010101001100101101",
"01000011010011110100110001000011",
"00010001001111010101001001001011",
"01001001010100100101010000000000",
"01010010010001010100011101000111",
"01000101010100100101000000101101",
"01001100010000010100001101010011",
"00111101010011110101001001000101",
"01010010010101000000000000001101",
"01000101010001110100011101001001",
"01001110010010010010110101010010",
"01010011010101000101010101010000",
"00101100001011010101001100011100",
"00000000000001010100001000001010",
"00000010010000000100011100001000",
"00001111000101100100110000000000",
"11001100010110000011111000001111",
"00100000000110010000111101010101",
"00000010111111111101000001000110",
"11111111110100000100011000100010",
"00001100001111010000100100000001",
"01000011010011110100110000000000",
"01001111010000110010110101001011",
"01000101010101000100111001010101",
"00011010000110100001101001010010",
"00011010000110100000111100100010",
"00010110111111111100000001000110",
"00010011001111010000100000000001",
"01010100010001010101001100000000",
"01010101010011110100001100101101",
"01010010010001010101010001001110",
"01010010010001010101001100101101",
"01000101010000110100100101010110",
"11000000010001100001101000011010",
"00111101000000100001011011111111",
"01000101010100110000000000001010",
"01010101010011110100001101010100",
"01010010010001010101010001001110",
"11111111110101000100011001000011",
"00001010011011001100011000000010",
"00000010000111011001000000010000",
"01010110000000101000100000010000",
"00010110000010101001000101010101",
"00100101000010101001000100010000",
"10001000000100001000100100010000",
"10001000000100000000000110010000",
"01000110000011100000000100011101",
"01000110000000011111111111011000",
"00110101000000100000101001010100",
"00000010000010101001100001000110",
"00100001010000100001110000101100",
"00001010011001000100011000000000",
"00000000001000000100011000000010",
"01000010000010100101101100101101",
"00001111010101010000000000000100",
"00100011010101000000101000100000",
"00000010000010100110100001000110",
"00000101010000100101101100010111",
"00111110010101110000111000000000",
"01010101000010001100101011110110",
"00000001000010101010010001000110",
"00000010000010101001110001000110",
"00000000000000110100001000101100",
"01000110111010101100000100111110",
"01000100000000011111111111010100",
"01010010000000000000101100111101",
"01000011010001000100000101000101",
"01010100010011100101010101001111",
"00000000000001100101001001000101",
"01000001010101000101001101010110",
"00000000000001110100101101000011",
"01001110010001010100110001010110",
"00000101010010000101010001000111",
"01000101010101110101001100000000",
"00000000000010000101000001000101",
"01000011010100110101100101010011",
"01001011010000110100111101001100",
"01001111010100110000000000001001",
"01000101010000110101001001010101",
"00000100010001000100100100101101",
"01101001011101000010001100000000",
"00111110000000000000001101100010",
"00000000000000110110111001101001",
"00000011011000100110100101110100",
"01000100010011000100100000000000",
"01000001010100000000000000000011",
"01001010000000000000100101000100",
"01010100010000010101011001000001",
"01010010010001010100110101001001",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000"
)
                           );
  type dvec is array (0 to 9 - 1) of DataVec;
  signal bdata: dvec;
  signal old: std_ulogic_vector(ROMrange'high downto 11);
  
begin
  
  fetch: process(Clock) is
  begin
    if rising_edge(Clock) then
         old <= Address(old'range);
	   for i in bdata'range loop
	     bData(i) <= ROM(i)(to_integer(std_ulogic_vector(Address(11 - 1 downto 2))) MOD blocks'length);
		end loop;
	 end if;
  end process fetch;

  Data <= 
          bdata(0 ) when unsigned(old) = 0 else
          bdata(1 ) when unsigned(old) = 1 else
          bdata(2 ) when unsigned(old) = 2 else
          bdata(3 ) when unsigned(old) = 3 else
          bdata(4 ) when unsigned(old) = 4 else
          bdata(5 ) when unsigned(old) = 5 else
          bdata(6 ) when unsigned(old) = 6 else
          bdata(7 ) when unsigned(old) = 7 else
          bdata(8 ) when unsigned(old) = 8 else
          (others => '0');
			 
end RTL;
